// ed_synth.v

// Generated using ACDS version 20.4 72

`timescale 1 ps / 1 ps
module ed_synth (
		input  wire       core_clk_iopll_reset_reset,               //             core_clk_iopll_reset.reset
		input  wire       core_clk_iopll_ref_clk_clk,               //           core_clk_iopll_ref_clk.clk
		input  wire       hbm_0_example_design_pll_ref_clk_clk,     // hbm_0_example_design_pll_ref_clk.clk
		input  wire       hbm_0_example_design_wmcrst_n_in_reset_n, // hbm_0_example_design_wmcrst_n_in.reset_n
		input  wire       hbm_only_reset_in_reset,                  //                hbm_only_reset_in.reset
		input  wire       m2u_bridge_cattrip,                       //                       m2u_bridge.cattrip
		input  wire [2:0] m2u_bridge_temp,                          //                                 .temp
		input  wire [7:0] m2u_bridge_wso,                           //                                 .wso
		output wire       m2u_bridge_reset_n,                       //                                 .reset_n
		output wire       m2u_bridge_wrst_n,                        //                                 .wrst_n
		output wire       m2u_bridge_wrck,                          //                                 .wrck
		output wire       m2u_bridge_shiftwr,                       //                                 .shiftwr
		output wire       m2u_bridge_capturewr,                     //                                 .capturewr
		output wire       m2u_bridge_updatewr,                      //                                 .updatewr
		output wire       m2u_bridge_selectwir,                     //                                 .selectwir
		output wire       m2u_bridge_wsi,                           //                                 .wsi
		output wire       tg0_0_status_traffic_gen_pass,            //                     tg0_0_status.traffic_gen_pass
		output wire       tg0_0_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg0_0_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg0_1_status_traffic_gen_pass,            //                     tg0_1_status.traffic_gen_pass
		output wire       tg0_1_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg0_1_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg1_0_status_traffic_gen_pass,            //                     tg1_0_status.traffic_gen_pass
		output wire       tg1_0_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg1_0_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg1_1_status_traffic_gen_pass,            //                     tg1_1_status.traffic_gen_pass
		output wire       tg1_1_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg1_1_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg2_0_status_traffic_gen_pass,            //                     tg2_0_status.traffic_gen_pass
		output wire       tg2_0_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg2_0_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg2_1_status_traffic_gen_pass,            //                     tg2_1_status.traffic_gen_pass
		output wire       tg2_1_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg2_1_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg3_0_status_traffic_gen_pass,            //                     tg3_0_status.traffic_gen_pass
		output wire       tg3_0_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg3_0_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg3_1_status_traffic_gen_pass,            //                     tg3_1_status.traffic_gen_pass
		output wire       tg3_1_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg3_1_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg4_0_status_traffic_gen_pass,            //                     tg4_0_status.traffic_gen_pass
		output wire       tg4_0_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg4_0_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg4_1_status_traffic_gen_pass,            //                     tg4_1_status.traffic_gen_pass
		output wire       tg4_1_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg4_1_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg5_0_status_traffic_gen_pass,            //                     tg5_0_status.traffic_gen_pass
		output wire       tg5_0_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg5_0_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg5_1_status_traffic_gen_pass,            //                     tg5_1_status.traffic_gen_pass
		output wire       tg5_1_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg5_1_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg6_0_status_traffic_gen_pass,            //                     tg6_0_status.traffic_gen_pass
		output wire       tg6_0_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg6_0_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg6_1_status_traffic_gen_pass,            //                     tg6_1_status.traffic_gen_pass
		output wire       tg6_1_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg6_1_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg7_0_status_traffic_gen_pass,            //                     tg7_0_status.traffic_gen_pass
		output wire       tg7_0_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg7_0_status_traffic_gen_timeout,         //                                 .traffic_gen_timeout
		output wire       tg7_1_status_traffic_gen_pass,            //                     tg7_1_status.traffic_gen_pass
		output wire       tg7_1_status_traffic_gen_fail,            //                                 .traffic_gen_fail
		output wire       tg7_1_status_traffic_gen_timeout          //                                 .traffic_gen_timeout
	);

	wire    [1:0] tg0_0_axi_awburst;                                // tg0_0:awburst -> hbm_0_example_design:axi_0_0_awburst
	wire    [0:0] tg0_0_axi_awuser;                                 // tg0_0:awuser_ap -> hbm_0_example_design:axi_0_0_awuser
	wire    [7:0] tg0_0_axi_arlen;                                  // tg0_0:arlen -> hbm_0_example_design:axi_0_0_arlen
	wire    [3:0] tg0_0_axi_arqos;                                  // tg0_0:arqos -> hbm_0_example_design:axi_0_0_arqos
	wire   [31:0] tg0_0_axi_wstrb;                                  // tg0_0:wstrb -> hbm_0_example_design:axi_0_0_wstrb
	wire          tg0_0_axi_wready;                                 // hbm_0_example_design:axi_0_0_wready -> tg0_0:wready
	wire    [6:0] tg0_0_axi_rid;                                    // hbm_0_example_design:axi_0_0_rid -> tg0_0:rid
	wire          tg0_0_axi_rready;                                 // tg0_0:rready -> hbm_0_example_design:axi_0_0_rready
	wire    [7:0] tg0_0_axi_awlen;                                  // tg0_0:awlen -> hbm_0_example_design:axi_0_0_awlen
	wire    [3:0] tg0_0_axi_awqos;                                  // tg0_0:awqos -> hbm_0_example_design:axi_0_0_awqos
	wire          tg0_0_axi_wvalid;                                 // tg0_0:wvalid -> hbm_0_example_design:axi_0_0_wvalid
	wire   [29:0] tg0_0_axi_araddr;                                 // tg0_0:araddr -> hbm_0_example_design:axi_0_0_araddr
	wire    [2:0] tg0_0_axi_arprot;                                 // tg0_0:arprot -> hbm_0_example_design:axi_0_0_arprot
	wire    [2:0] tg0_0_axi_awprot;                                 // tg0_0:awprot -> hbm_0_example_design:axi_0_0_awprot
	wire  [255:0] tg0_0_axi_wdata;                                  // tg0_0:wdata -> hbm_0_example_design:axi_0_0_wdata
	wire          tg0_0_axi_arvalid;                                // tg0_0:arvalid -> hbm_0_example_design:axi_0_0_arvalid
	wire    [6:0] tg0_0_axi_arid;                                   // tg0_0:arid -> hbm_0_example_design:axi_0_0_arid
	wire   [29:0] tg0_0_axi_awaddr;                                 // tg0_0:awaddr -> hbm_0_example_design:axi_0_0_awaddr
	wire    [1:0] tg0_0_axi_bresp;                                  // hbm_0_example_design:axi_0_0_bresp -> tg0_0:bresp
	wire          tg0_0_axi_arready;                                // hbm_0_example_design:axi_0_0_arready -> tg0_0:arready
	wire  [255:0] tg0_0_axi_rdata;                                  // hbm_0_example_design:axi_0_0_rdata -> tg0_0:rdata
	wire          tg0_0_axi_awready;                                // hbm_0_example_design:axi_0_0_awready -> tg0_0:awready
	wire    [1:0] tg0_0_axi_arburst;                                // tg0_0:arburst -> hbm_0_example_design:axi_0_0_arburst
	wire    [2:0] tg0_0_axi_arsize;                                 // tg0_0:arsize -> hbm_0_example_design:axi_0_0_arsize
	wire          tg0_0_axi_bready;                                 // tg0_0:bready -> hbm_0_example_design:axi_0_0_bready
	wire          tg0_0_axi_rlast;                                  // hbm_0_example_design:axi_0_0_rlast -> tg0_0:rlast
	wire          tg0_0_axi_wlast;                                  // tg0_0:wlast -> hbm_0_example_design:axi_0_0_wlast
	wire    [1:0] tg0_0_axi_rresp;                                  // hbm_0_example_design:axi_0_0_rresp -> tg0_0:rresp
	wire    [6:0] tg0_0_axi_awid;                                   // tg0_0:awid -> hbm_0_example_design:axi_0_0_awid
	wire    [6:0] tg0_0_axi_bid;                                    // hbm_0_example_design:axi_0_0_bid -> tg0_0:bid
	wire          tg0_0_axi_bvalid;                                 // hbm_0_example_design:axi_0_0_bvalid -> tg0_0:bvalid
	wire    [2:0] tg0_0_axi_awsize;                                 // tg0_0:awsize -> hbm_0_example_design:axi_0_0_awsize
	wire          tg0_0_axi_awvalid;                                // tg0_0:awvalid -> hbm_0_example_design:axi_0_0_awvalid
	wire    [0:0] tg0_0_axi_aruser;                                 // tg0_0:aruser_ap -> hbm_0_example_design:axi_0_0_aruser
	wire          tg0_0_axi_rvalid;                                 // hbm_0_example_design:axi_0_0_rvalid -> tg0_0:rvalid
	wire    [1:0] tg0_1_axi_awburst;                                // tg0_1:awburst -> hbm_0_example_design:axi_0_1_awburst
	wire    [0:0] tg0_1_axi_awuser;                                 // tg0_1:awuser_ap -> hbm_0_example_design:axi_0_1_awuser
	wire    [7:0] tg0_1_axi_arlen;                                  // tg0_1:arlen -> hbm_0_example_design:axi_0_1_arlen
	wire    [3:0] tg0_1_axi_arqos;                                  // tg0_1:arqos -> hbm_0_example_design:axi_0_1_arqos
	wire   [31:0] tg0_1_axi_wstrb;                                  // tg0_1:wstrb -> hbm_0_example_design:axi_0_1_wstrb
	wire          tg0_1_axi_wready;                                 // hbm_0_example_design:axi_0_1_wready -> tg0_1:wready
	wire    [6:0] tg0_1_axi_rid;                                    // hbm_0_example_design:axi_0_1_rid -> tg0_1:rid
	wire          tg0_1_axi_rready;                                 // tg0_1:rready -> hbm_0_example_design:axi_0_1_rready
	wire    [7:0] tg0_1_axi_awlen;                                  // tg0_1:awlen -> hbm_0_example_design:axi_0_1_awlen
	wire    [3:0] tg0_1_axi_awqos;                                  // tg0_1:awqos -> hbm_0_example_design:axi_0_1_awqos
	wire          tg0_1_axi_wvalid;                                 // tg0_1:wvalid -> hbm_0_example_design:axi_0_1_wvalid
	wire   [29:0] tg0_1_axi_araddr;                                 // tg0_1:araddr -> hbm_0_example_design:axi_0_1_araddr
	wire    [2:0] tg0_1_axi_arprot;                                 // tg0_1:arprot -> hbm_0_example_design:axi_0_1_arprot
	wire    [2:0] tg0_1_axi_awprot;                                 // tg0_1:awprot -> hbm_0_example_design:axi_0_1_awprot
	wire  [255:0] tg0_1_axi_wdata;                                  // tg0_1:wdata -> hbm_0_example_design:axi_0_1_wdata
	wire          tg0_1_axi_arvalid;                                // tg0_1:arvalid -> hbm_0_example_design:axi_0_1_arvalid
	wire    [6:0] tg0_1_axi_arid;                                   // tg0_1:arid -> hbm_0_example_design:axi_0_1_arid
	wire   [29:0] tg0_1_axi_awaddr;                                 // tg0_1:awaddr -> hbm_0_example_design:axi_0_1_awaddr
	wire    [1:0] tg0_1_axi_bresp;                                  // hbm_0_example_design:axi_0_1_bresp -> tg0_1:bresp
	wire          tg0_1_axi_arready;                                // hbm_0_example_design:axi_0_1_arready -> tg0_1:arready
	wire  [255:0] tg0_1_axi_rdata;                                  // hbm_0_example_design:axi_0_1_rdata -> tg0_1:rdata
	wire          tg0_1_axi_awready;                                // hbm_0_example_design:axi_0_1_awready -> tg0_1:awready
	wire    [1:0] tg0_1_axi_arburst;                                // tg0_1:arburst -> hbm_0_example_design:axi_0_1_arburst
	wire    [2:0] tg0_1_axi_arsize;                                 // tg0_1:arsize -> hbm_0_example_design:axi_0_1_arsize
	wire          tg0_1_axi_bready;                                 // tg0_1:bready -> hbm_0_example_design:axi_0_1_bready
	wire          tg0_1_axi_rlast;                                  // hbm_0_example_design:axi_0_1_rlast -> tg0_1:rlast
	wire          tg0_1_axi_wlast;                                  // tg0_1:wlast -> hbm_0_example_design:axi_0_1_wlast
	wire    [1:0] tg0_1_axi_rresp;                                  // hbm_0_example_design:axi_0_1_rresp -> tg0_1:rresp
	wire    [6:0] tg0_1_axi_awid;                                   // tg0_1:awid -> hbm_0_example_design:axi_0_1_awid
	wire    [6:0] tg0_1_axi_bid;                                    // hbm_0_example_design:axi_0_1_bid -> tg0_1:bid
	wire          tg0_1_axi_bvalid;                                 // hbm_0_example_design:axi_0_1_bvalid -> tg0_1:bvalid
	wire    [2:0] tg0_1_axi_awsize;                                 // tg0_1:awsize -> hbm_0_example_design:axi_0_1_awsize
	wire          tg0_1_axi_awvalid;                                // tg0_1:awvalid -> hbm_0_example_design:axi_0_1_awvalid
	wire    [0:0] tg0_1_axi_aruser;                                 // tg0_1:aruser_ap -> hbm_0_example_design:axi_0_1_aruser
	wire          tg0_1_axi_rvalid;                                 // hbm_0_example_design:axi_0_1_rvalid -> tg0_1:rvalid
	wire    [1:0] tg1_0_axi_awburst;                                // tg1_0:awburst -> hbm_0_example_design:axi_1_0_awburst
	wire    [0:0] tg1_0_axi_awuser;                                 // tg1_0:awuser_ap -> hbm_0_example_design:axi_1_0_awuser
	wire    [7:0] tg1_0_axi_arlen;                                  // tg1_0:arlen -> hbm_0_example_design:axi_1_0_arlen
	wire    [3:0] tg1_0_axi_arqos;                                  // tg1_0:arqos -> hbm_0_example_design:axi_1_0_arqos
	wire   [31:0] tg1_0_axi_wstrb;                                  // tg1_0:wstrb -> hbm_0_example_design:axi_1_0_wstrb
	wire          tg1_0_axi_wready;                                 // hbm_0_example_design:axi_1_0_wready -> tg1_0:wready
	wire    [6:0] tg1_0_axi_rid;                                    // hbm_0_example_design:axi_1_0_rid -> tg1_0:rid
	wire          tg1_0_axi_rready;                                 // tg1_0:rready -> hbm_0_example_design:axi_1_0_rready
	wire    [7:0] tg1_0_axi_awlen;                                  // tg1_0:awlen -> hbm_0_example_design:axi_1_0_awlen
	wire    [3:0] tg1_0_axi_awqos;                                  // tg1_0:awqos -> hbm_0_example_design:axi_1_0_awqos
	wire          tg1_0_axi_wvalid;                                 // tg1_0:wvalid -> hbm_0_example_design:axi_1_0_wvalid
	wire   [29:0] tg1_0_axi_araddr;                                 // tg1_0:araddr -> hbm_0_example_design:axi_1_0_araddr
	wire    [2:0] tg1_0_axi_arprot;                                 // tg1_0:arprot -> hbm_0_example_design:axi_1_0_arprot
	wire    [2:0] tg1_0_axi_awprot;                                 // tg1_0:awprot -> hbm_0_example_design:axi_1_0_awprot
	wire  [255:0] tg1_0_axi_wdata;                                  // tg1_0:wdata -> hbm_0_example_design:axi_1_0_wdata
	wire          tg1_0_axi_arvalid;                                // tg1_0:arvalid -> hbm_0_example_design:axi_1_0_arvalid
	wire    [6:0] tg1_0_axi_arid;                                   // tg1_0:arid -> hbm_0_example_design:axi_1_0_arid
	wire   [29:0] tg1_0_axi_awaddr;                                 // tg1_0:awaddr -> hbm_0_example_design:axi_1_0_awaddr
	wire    [1:0] tg1_0_axi_bresp;                                  // hbm_0_example_design:axi_1_0_bresp -> tg1_0:bresp
	wire          tg1_0_axi_arready;                                // hbm_0_example_design:axi_1_0_arready -> tg1_0:arready
	wire  [255:0] tg1_0_axi_rdata;                                  // hbm_0_example_design:axi_1_0_rdata -> tg1_0:rdata
	wire          tg1_0_axi_awready;                                // hbm_0_example_design:axi_1_0_awready -> tg1_0:awready
	wire    [1:0] tg1_0_axi_arburst;                                // tg1_0:arburst -> hbm_0_example_design:axi_1_0_arburst
	wire    [2:0] tg1_0_axi_arsize;                                 // tg1_0:arsize -> hbm_0_example_design:axi_1_0_arsize
	wire          tg1_0_axi_bready;                                 // tg1_0:bready -> hbm_0_example_design:axi_1_0_bready
	wire          tg1_0_axi_rlast;                                  // hbm_0_example_design:axi_1_0_rlast -> tg1_0:rlast
	wire          tg1_0_axi_wlast;                                  // tg1_0:wlast -> hbm_0_example_design:axi_1_0_wlast
	wire    [1:0] tg1_0_axi_rresp;                                  // hbm_0_example_design:axi_1_0_rresp -> tg1_0:rresp
	wire    [6:0] tg1_0_axi_awid;                                   // tg1_0:awid -> hbm_0_example_design:axi_1_0_awid
	wire    [6:0] tg1_0_axi_bid;                                    // hbm_0_example_design:axi_1_0_bid -> tg1_0:bid
	wire          tg1_0_axi_bvalid;                                 // hbm_0_example_design:axi_1_0_bvalid -> tg1_0:bvalid
	wire    [2:0] tg1_0_axi_awsize;                                 // tg1_0:awsize -> hbm_0_example_design:axi_1_0_awsize
	wire          tg1_0_axi_awvalid;                                // tg1_0:awvalid -> hbm_0_example_design:axi_1_0_awvalid
	wire    [0:0] tg1_0_axi_aruser;                                 // tg1_0:aruser_ap -> hbm_0_example_design:axi_1_0_aruser
	wire          tg1_0_axi_rvalid;                                 // hbm_0_example_design:axi_1_0_rvalid -> tg1_0:rvalid
	wire    [1:0] tg1_1_axi_awburst;                                // tg1_1:awburst -> hbm_0_example_design:axi_1_1_awburst
	wire    [0:0] tg1_1_axi_awuser;                                 // tg1_1:awuser_ap -> hbm_0_example_design:axi_1_1_awuser
	wire    [7:0] tg1_1_axi_arlen;                                  // tg1_1:arlen -> hbm_0_example_design:axi_1_1_arlen
	wire    [3:0] tg1_1_axi_arqos;                                  // tg1_1:arqos -> hbm_0_example_design:axi_1_1_arqos
	wire   [31:0] tg1_1_axi_wstrb;                                  // tg1_1:wstrb -> hbm_0_example_design:axi_1_1_wstrb
	wire          tg1_1_axi_wready;                                 // hbm_0_example_design:axi_1_1_wready -> tg1_1:wready
	wire    [6:0] tg1_1_axi_rid;                                    // hbm_0_example_design:axi_1_1_rid -> tg1_1:rid
	wire          tg1_1_axi_rready;                                 // tg1_1:rready -> hbm_0_example_design:axi_1_1_rready
	wire    [7:0] tg1_1_axi_awlen;                                  // tg1_1:awlen -> hbm_0_example_design:axi_1_1_awlen
	wire    [3:0] tg1_1_axi_awqos;                                  // tg1_1:awqos -> hbm_0_example_design:axi_1_1_awqos
	wire          tg1_1_axi_wvalid;                                 // tg1_1:wvalid -> hbm_0_example_design:axi_1_1_wvalid
	wire   [29:0] tg1_1_axi_araddr;                                 // tg1_1:araddr -> hbm_0_example_design:axi_1_1_araddr
	wire    [2:0] tg1_1_axi_arprot;                                 // tg1_1:arprot -> hbm_0_example_design:axi_1_1_arprot
	wire    [2:0] tg1_1_axi_awprot;                                 // tg1_1:awprot -> hbm_0_example_design:axi_1_1_awprot
	wire  [255:0] tg1_1_axi_wdata;                                  // tg1_1:wdata -> hbm_0_example_design:axi_1_1_wdata
	wire          tg1_1_axi_arvalid;                                // tg1_1:arvalid -> hbm_0_example_design:axi_1_1_arvalid
	wire    [6:0] tg1_1_axi_arid;                                   // tg1_1:arid -> hbm_0_example_design:axi_1_1_arid
	wire   [29:0] tg1_1_axi_awaddr;                                 // tg1_1:awaddr -> hbm_0_example_design:axi_1_1_awaddr
	wire    [1:0] tg1_1_axi_bresp;                                  // hbm_0_example_design:axi_1_1_bresp -> tg1_1:bresp
	wire          tg1_1_axi_arready;                                // hbm_0_example_design:axi_1_1_arready -> tg1_1:arready
	wire  [255:0] tg1_1_axi_rdata;                                  // hbm_0_example_design:axi_1_1_rdata -> tg1_1:rdata
	wire          tg1_1_axi_awready;                                // hbm_0_example_design:axi_1_1_awready -> tg1_1:awready
	wire    [1:0] tg1_1_axi_arburst;                                // tg1_1:arburst -> hbm_0_example_design:axi_1_1_arburst
	wire    [2:0] tg1_1_axi_arsize;                                 // tg1_1:arsize -> hbm_0_example_design:axi_1_1_arsize
	wire          tg1_1_axi_bready;                                 // tg1_1:bready -> hbm_0_example_design:axi_1_1_bready
	wire          tg1_1_axi_rlast;                                  // hbm_0_example_design:axi_1_1_rlast -> tg1_1:rlast
	wire          tg1_1_axi_wlast;                                  // tg1_1:wlast -> hbm_0_example_design:axi_1_1_wlast
	wire    [1:0] tg1_1_axi_rresp;                                  // hbm_0_example_design:axi_1_1_rresp -> tg1_1:rresp
	wire    [6:0] tg1_1_axi_awid;                                   // tg1_1:awid -> hbm_0_example_design:axi_1_1_awid
	wire    [6:0] tg1_1_axi_bid;                                    // hbm_0_example_design:axi_1_1_bid -> tg1_1:bid
	wire          tg1_1_axi_bvalid;                                 // hbm_0_example_design:axi_1_1_bvalid -> tg1_1:bvalid
	wire    [2:0] tg1_1_axi_awsize;                                 // tg1_1:awsize -> hbm_0_example_design:axi_1_1_awsize
	wire          tg1_1_axi_awvalid;                                // tg1_1:awvalid -> hbm_0_example_design:axi_1_1_awvalid
	wire    [0:0] tg1_1_axi_aruser;                                 // tg1_1:aruser_ap -> hbm_0_example_design:axi_1_1_aruser
	wire          tg1_1_axi_rvalid;                                 // hbm_0_example_design:axi_1_1_rvalid -> tg1_1:rvalid
	wire    [1:0] tg2_0_axi_awburst;                                // tg2_0:awburst -> hbm_0_example_design:axi_2_0_awburst
	wire    [0:0] tg2_0_axi_awuser;                                 // tg2_0:awuser_ap -> hbm_0_example_design:axi_2_0_awuser
	wire    [7:0] tg2_0_axi_arlen;                                  // tg2_0:arlen -> hbm_0_example_design:axi_2_0_arlen
	wire    [3:0] tg2_0_axi_arqos;                                  // tg2_0:arqos -> hbm_0_example_design:axi_2_0_arqos
	wire   [31:0] tg2_0_axi_wstrb;                                  // tg2_0:wstrb -> hbm_0_example_design:axi_2_0_wstrb
	wire          tg2_0_axi_wready;                                 // hbm_0_example_design:axi_2_0_wready -> tg2_0:wready
	wire    [6:0] tg2_0_axi_rid;                                    // hbm_0_example_design:axi_2_0_rid -> tg2_0:rid
	wire          tg2_0_axi_rready;                                 // tg2_0:rready -> hbm_0_example_design:axi_2_0_rready
	wire    [7:0] tg2_0_axi_awlen;                                  // tg2_0:awlen -> hbm_0_example_design:axi_2_0_awlen
	wire    [3:0] tg2_0_axi_awqos;                                  // tg2_0:awqos -> hbm_0_example_design:axi_2_0_awqos
	wire          tg2_0_axi_wvalid;                                 // tg2_0:wvalid -> hbm_0_example_design:axi_2_0_wvalid
	wire   [29:0] tg2_0_axi_araddr;                                 // tg2_0:araddr -> hbm_0_example_design:axi_2_0_araddr
	wire    [2:0] tg2_0_axi_arprot;                                 // tg2_0:arprot -> hbm_0_example_design:axi_2_0_arprot
	wire    [2:0] tg2_0_axi_awprot;                                 // tg2_0:awprot -> hbm_0_example_design:axi_2_0_awprot
	wire  [255:0] tg2_0_axi_wdata;                                  // tg2_0:wdata -> hbm_0_example_design:axi_2_0_wdata
	wire          tg2_0_axi_arvalid;                                // tg2_0:arvalid -> hbm_0_example_design:axi_2_0_arvalid
	wire    [6:0] tg2_0_axi_arid;                                   // tg2_0:arid -> hbm_0_example_design:axi_2_0_arid
	wire   [29:0] tg2_0_axi_awaddr;                                 // tg2_0:awaddr -> hbm_0_example_design:axi_2_0_awaddr
	wire    [1:0] tg2_0_axi_bresp;                                  // hbm_0_example_design:axi_2_0_bresp -> tg2_0:bresp
	wire          tg2_0_axi_arready;                                // hbm_0_example_design:axi_2_0_arready -> tg2_0:arready
	wire  [255:0] tg2_0_axi_rdata;                                  // hbm_0_example_design:axi_2_0_rdata -> tg2_0:rdata
	wire          tg2_0_axi_awready;                                // hbm_0_example_design:axi_2_0_awready -> tg2_0:awready
	wire    [1:0] tg2_0_axi_arburst;                                // tg2_0:arburst -> hbm_0_example_design:axi_2_0_arburst
	wire    [2:0] tg2_0_axi_arsize;                                 // tg2_0:arsize -> hbm_0_example_design:axi_2_0_arsize
	wire          tg2_0_axi_bready;                                 // tg2_0:bready -> hbm_0_example_design:axi_2_0_bready
	wire          tg2_0_axi_rlast;                                  // hbm_0_example_design:axi_2_0_rlast -> tg2_0:rlast
	wire          tg2_0_axi_wlast;                                  // tg2_0:wlast -> hbm_0_example_design:axi_2_0_wlast
	wire    [1:0] tg2_0_axi_rresp;                                  // hbm_0_example_design:axi_2_0_rresp -> tg2_0:rresp
	wire    [6:0] tg2_0_axi_awid;                                   // tg2_0:awid -> hbm_0_example_design:axi_2_0_awid
	wire    [6:0] tg2_0_axi_bid;                                    // hbm_0_example_design:axi_2_0_bid -> tg2_0:bid
	wire          tg2_0_axi_bvalid;                                 // hbm_0_example_design:axi_2_0_bvalid -> tg2_0:bvalid
	wire    [2:0] tg2_0_axi_awsize;                                 // tg2_0:awsize -> hbm_0_example_design:axi_2_0_awsize
	wire          tg2_0_axi_awvalid;                                // tg2_0:awvalid -> hbm_0_example_design:axi_2_0_awvalid
	wire    [0:0] tg2_0_axi_aruser;                                 // tg2_0:aruser_ap -> hbm_0_example_design:axi_2_0_aruser
	wire          tg2_0_axi_rvalid;                                 // hbm_0_example_design:axi_2_0_rvalid -> tg2_0:rvalid
	wire    [1:0] tg2_1_axi_awburst;                                // tg2_1:awburst -> hbm_0_example_design:axi_2_1_awburst
	wire    [0:0] tg2_1_axi_awuser;                                 // tg2_1:awuser_ap -> hbm_0_example_design:axi_2_1_awuser
	wire    [7:0] tg2_1_axi_arlen;                                  // tg2_1:arlen -> hbm_0_example_design:axi_2_1_arlen
	wire    [3:0] tg2_1_axi_arqos;                                  // tg2_1:arqos -> hbm_0_example_design:axi_2_1_arqos
	wire   [31:0] tg2_1_axi_wstrb;                                  // tg2_1:wstrb -> hbm_0_example_design:axi_2_1_wstrb
	wire          tg2_1_axi_wready;                                 // hbm_0_example_design:axi_2_1_wready -> tg2_1:wready
	wire    [6:0] tg2_1_axi_rid;                                    // hbm_0_example_design:axi_2_1_rid -> tg2_1:rid
	wire          tg2_1_axi_rready;                                 // tg2_1:rready -> hbm_0_example_design:axi_2_1_rready
	wire    [7:0] tg2_1_axi_awlen;                                  // tg2_1:awlen -> hbm_0_example_design:axi_2_1_awlen
	wire    [3:0] tg2_1_axi_awqos;                                  // tg2_1:awqos -> hbm_0_example_design:axi_2_1_awqos
	wire          tg2_1_axi_wvalid;                                 // tg2_1:wvalid -> hbm_0_example_design:axi_2_1_wvalid
	wire   [29:0] tg2_1_axi_araddr;                                 // tg2_1:araddr -> hbm_0_example_design:axi_2_1_araddr
	wire    [2:0] tg2_1_axi_arprot;                                 // tg2_1:arprot -> hbm_0_example_design:axi_2_1_arprot
	wire    [2:0] tg2_1_axi_awprot;                                 // tg2_1:awprot -> hbm_0_example_design:axi_2_1_awprot
	wire  [255:0] tg2_1_axi_wdata;                                  // tg2_1:wdata -> hbm_0_example_design:axi_2_1_wdata
	wire          tg2_1_axi_arvalid;                                // tg2_1:arvalid -> hbm_0_example_design:axi_2_1_arvalid
	wire    [6:0] tg2_1_axi_arid;                                   // tg2_1:arid -> hbm_0_example_design:axi_2_1_arid
	wire   [29:0] tg2_1_axi_awaddr;                                 // tg2_1:awaddr -> hbm_0_example_design:axi_2_1_awaddr
	wire    [1:0] tg2_1_axi_bresp;                                  // hbm_0_example_design:axi_2_1_bresp -> tg2_1:bresp
	wire          tg2_1_axi_arready;                                // hbm_0_example_design:axi_2_1_arready -> tg2_1:arready
	wire  [255:0] tg2_1_axi_rdata;                                  // hbm_0_example_design:axi_2_1_rdata -> tg2_1:rdata
	wire          tg2_1_axi_awready;                                // hbm_0_example_design:axi_2_1_awready -> tg2_1:awready
	wire    [1:0] tg2_1_axi_arburst;                                // tg2_1:arburst -> hbm_0_example_design:axi_2_1_arburst
	wire    [2:0] tg2_1_axi_arsize;                                 // tg2_1:arsize -> hbm_0_example_design:axi_2_1_arsize
	wire          tg2_1_axi_bready;                                 // tg2_1:bready -> hbm_0_example_design:axi_2_1_bready
	wire          tg2_1_axi_rlast;                                  // hbm_0_example_design:axi_2_1_rlast -> tg2_1:rlast
	wire          tg2_1_axi_wlast;                                  // tg2_1:wlast -> hbm_0_example_design:axi_2_1_wlast
	wire    [1:0] tg2_1_axi_rresp;                                  // hbm_0_example_design:axi_2_1_rresp -> tg2_1:rresp
	wire    [6:0] tg2_1_axi_awid;                                   // tg2_1:awid -> hbm_0_example_design:axi_2_1_awid
	wire    [6:0] tg2_1_axi_bid;                                    // hbm_0_example_design:axi_2_1_bid -> tg2_1:bid
	wire          tg2_1_axi_bvalid;                                 // hbm_0_example_design:axi_2_1_bvalid -> tg2_1:bvalid
	wire    [2:0] tg2_1_axi_awsize;                                 // tg2_1:awsize -> hbm_0_example_design:axi_2_1_awsize
	wire          tg2_1_axi_awvalid;                                // tg2_1:awvalid -> hbm_0_example_design:axi_2_1_awvalid
	wire    [0:0] tg2_1_axi_aruser;                                 // tg2_1:aruser_ap -> hbm_0_example_design:axi_2_1_aruser
	wire          tg2_1_axi_rvalid;                                 // hbm_0_example_design:axi_2_1_rvalid -> tg2_1:rvalid
	wire    [1:0] tg3_0_axi_awburst;                                // tg3_0:awburst -> hbm_0_example_design:axi_3_0_awburst
	wire    [0:0] tg3_0_axi_awuser;                                 // tg3_0:awuser_ap -> hbm_0_example_design:axi_3_0_awuser
	wire    [7:0] tg3_0_axi_arlen;                                  // tg3_0:arlen -> hbm_0_example_design:axi_3_0_arlen
	wire    [3:0] tg3_0_axi_arqos;                                  // tg3_0:arqos -> hbm_0_example_design:axi_3_0_arqos
	wire   [31:0] tg3_0_axi_wstrb;                                  // tg3_0:wstrb -> hbm_0_example_design:axi_3_0_wstrb
	wire          tg3_0_axi_wready;                                 // hbm_0_example_design:axi_3_0_wready -> tg3_0:wready
	wire    [6:0] tg3_0_axi_rid;                                    // hbm_0_example_design:axi_3_0_rid -> tg3_0:rid
	wire          tg3_0_axi_rready;                                 // tg3_0:rready -> hbm_0_example_design:axi_3_0_rready
	wire    [7:0] tg3_0_axi_awlen;                                  // tg3_0:awlen -> hbm_0_example_design:axi_3_0_awlen
	wire    [3:0] tg3_0_axi_awqos;                                  // tg3_0:awqos -> hbm_0_example_design:axi_3_0_awqos
	wire          tg3_0_axi_wvalid;                                 // tg3_0:wvalid -> hbm_0_example_design:axi_3_0_wvalid
	wire   [29:0] tg3_0_axi_araddr;                                 // tg3_0:araddr -> hbm_0_example_design:axi_3_0_araddr
	wire    [2:0] tg3_0_axi_arprot;                                 // tg3_0:arprot -> hbm_0_example_design:axi_3_0_arprot
	wire    [2:0] tg3_0_axi_awprot;                                 // tg3_0:awprot -> hbm_0_example_design:axi_3_0_awprot
	wire  [255:0] tg3_0_axi_wdata;                                  // tg3_0:wdata -> hbm_0_example_design:axi_3_0_wdata
	wire          tg3_0_axi_arvalid;                                // tg3_0:arvalid -> hbm_0_example_design:axi_3_0_arvalid
	wire    [6:0] tg3_0_axi_arid;                                   // tg3_0:arid -> hbm_0_example_design:axi_3_0_arid
	wire   [29:0] tg3_0_axi_awaddr;                                 // tg3_0:awaddr -> hbm_0_example_design:axi_3_0_awaddr
	wire    [1:0] tg3_0_axi_bresp;                                  // hbm_0_example_design:axi_3_0_bresp -> tg3_0:bresp
	wire          tg3_0_axi_arready;                                // hbm_0_example_design:axi_3_0_arready -> tg3_0:arready
	wire  [255:0] tg3_0_axi_rdata;                                  // hbm_0_example_design:axi_3_0_rdata -> tg3_0:rdata
	wire          tg3_0_axi_awready;                                // hbm_0_example_design:axi_3_0_awready -> tg3_0:awready
	wire    [1:0] tg3_0_axi_arburst;                                // tg3_0:arburst -> hbm_0_example_design:axi_3_0_arburst
	wire    [2:0] tg3_0_axi_arsize;                                 // tg3_0:arsize -> hbm_0_example_design:axi_3_0_arsize
	wire          tg3_0_axi_bready;                                 // tg3_0:bready -> hbm_0_example_design:axi_3_0_bready
	wire          tg3_0_axi_rlast;                                  // hbm_0_example_design:axi_3_0_rlast -> tg3_0:rlast
	wire          tg3_0_axi_wlast;                                  // tg3_0:wlast -> hbm_0_example_design:axi_3_0_wlast
	wire    [1:0] tg3_0_axi_rresp;                                  // hbm_0_example_design:axi_3_0_rresp -> tg3_0:rresp
	wire    [6:0] tg3_0_axi_awid;                                   // tg3_0:awid -> hbm_0_example_design:axi_3_0_awid
	wire    [6:0] tg3_0_axi_bid;                                    // hbm_0_example_design:axi_3_0_bid -> tg3_0:bid
	wire          tg3_0_axi_bvalid;                                 // hbm_0_example_design:axi_3_0_bvalid -> tg3_0:bvalid
	wire    [2:0] tg3_0_axi_awsize;                                 // tg3_0:awsize -> hbm_0_example_design:axi_3_0_awsize
	wire          tg3_0_axi_awvalid;                                // tg3_0:awvalid -> hbm_0_example_design:axi_3_0_awvalid
	wire    [0:0] tg3_0_axi_aruser;                                 // tg3_0:aruser_ap -> hbm_0_example_design:axi_3_0_aruser
	wire          tg3_0_axi_rvalid;                                 // hbm_0_example_design:axi_3_0_rvalid -> tg3_0:rvalid
	wire    [1:0] tg3_1_axi_awburst;                                // tg3_1:awburst -> hbm_0_example_design:axi_3_1_awburst
	wire    [0:0] tg3_1_axi_awuser;                                 // tg3_1:awuser_ap -> hbm_0_example_design:axi_3_1_awuser
	wire    [7:0] tg3_1_axi_arlen;                                  // tg3_1:arlen -> hbm_0_example_design:axi_3_1_arlen
	wire    [3:0] tg3_1_axi_arqos;                                  // tg3_1:arqos -> hbm_0_example_design:axi_3_1_arqos
	wire   [31:0] tg3_1_axi_wstrb;                                  // tg3_1:wstrb -> hbm_0_example_design:axi_3_1_wstrb
	wire          tg3_1_axi_wready;                                 // hbm_0_example_design:axi_3_1_wready -> tg3_1:wready
	wire    [6:0] tg3_1_axi_rid;                                    // hbm_0_example_design:axi_3_1_rid -> tg3_1:rid
	wire          tg3_1_axi_rready;                                 // tg3_1:rready -> hbm_0_example_design:axi_3_1_rready
	wire    [7:0] tg3_1_axi_awlen;                                  // tg3_1:awlen -> hbm_0_example_design:axi_3_1_awlen
	wire    [3:0] tg3_1_axi_awqos;                                  // tg3_1:awqos -> hbm_0_example_design:axi_3_1_awqos
	wire          tg3_1_axi_wvalid;                                 // tg3_1:wvalid -> hbm_0_example_design:axi_3_1_wvalid
	wire   [29:0] tg3_1_axi_araddr;                                 // tg3_1:araddr -> hbm_0_example_design:axi_3_1_araddr
	wire    [2:0] tg3_1_axi_arprot;                                 // tg3_1:arprot -> hbm_0_example_design:axi_3_1_arprot
	wire    [2:0] tg3_1_axi_awprot;                                 // tg3_1:awprot -> hbm_0_example_design:axi_3_1_awprot
	wire  [255:0] tg3_1_axi_wdata;                                  // tg3_1:wdata -> hbm_0_example_design:axi_3_1_wdata
	wire          tg3_1_axi_arvalid;                                // tg3_1:arvalid -> hbm_0_example_design:axi_3_1_arvalid
	wire    [6:0] tg3_1_axi_arid;                                   // tg3_1:arid -> hbm_0_example_design:axi_3_1_arid
	wire   [29:0] tg3_1_axi_awaddr;                                 // tg3_1:awaddr -> hbm_0_example_design:axi_3_1_awaddr
	wire    [1:0] tg3_1_axi_bresp;                                  // hbm_0_example_design:axi_3_1_bresp -> tg3_1:bresp
	wire          tg3_1_axi_arready;                                // hbm_0_example_design:axi_3_1_arready -> tg3_1:arready
	wire  [255:0] tg3_1_axi_rdata;                                  // hbm_0_example_design:axi_3_1_rdata -> tg3_1:rdata
	wire          tg3_1_axi_awready;                                // hbm_0_example_design:axi_3_1_awready -> tg3_1:awready
	wire    [1:0] tg3_1_axi_arburst;                                // tg3_1:arburst -> hbm_0_example_design:axi_3_1_arburst
	wire    [2:0] tg3_1_axi_arsize;                                 // tg3_1:arsize -> hbm_0_example_design:axi_3_1_arsize
	wire          tg3_1_axi_bready;                                 // tg3_1:bready -> hbm_0_example_design:axi_3_1_bready
	wire          tg3_1_axi_rlast;                                  // hbm_0_example_design:axi_3_1_rlast -> tg3_1:rlast
	wire          tg3_1_axi_wlast;                                  // tg3_1:wlast -> hbm_0_example_design:axi_3_1_wlast
	wire    [1:0] tg3_1_axi_rresp;                                  // hbm_0_example_design:axi_3_1_rresp -> tg3_1:rresp
	wire    [6:0] tg3_1_axi_awid;                                   // tg3_1:awid -> hbm_0_example_design:axi_3_1_awid
	wire    [6:0] tg3_1_axi_bid;                                    // hbm_0_example_design:axi_3_1_bid -> tg3_1:bid
	wire          tg3_1_axi_bvalid;                                 // hbm_0_example_design:axi_3_1_bvalid -> tg3_1:bvalid
	wire    [2:0] tg3_1_axi_awsize;                                 // tg3_1:awsize -> hbm_0_example_design:axi_3_1_awsize
	wire          tg3_1_axi_awvalid;                                // tg3_1:awvalid -> hbm_0_example_design:axi_3_1_awvalid
	wire    [0:0] tg3_1_axi_aruser;                                 // tg3_1:aruser_ap -> hbm_0_example_design:axi_3_1_aruser
	wire          tg3_1_axi_rvalid;                                 // hbm_0_example_design:axi_3_1_rvalid -> tg3_1:rvalid
	wire    [1:0] tg4_0_axi_awburst;                                // tg4_0:awburst -> hbm_0_example_design:axi_4_0_awburst
	wire    [0:0] tg4_0_axi_awuser;                                 // tg4_0:awuser_ap -> hbm_0_example_design:axi_4_0_awuser
	wire    [7:0] tg4_0_axi_arlen;                                  // tg4_0:arlen -> hbm_0_example_design:axi_4_0_arlen
	wire    [3:0] tg4_0_axi_arqos;                                  // tg4_0:arqos -> hbm_0_example_design:axi_4_0_arqos
	wire   [31:0] tg4_0_axi_wstrb;                                  // tg4_0:wstrb -> hbm_0_example_design:axi_4_0_wstrb
	wire          tg4_0_axi_wready;                                 // hbm_0_example_design:axi_4_0_wready -> tg4_0:wready
	wire    [6:0] tg4_0_axi_rid;                                    // hbm_0_example_design:axi_4_0_rid -> tg4_0:rid
	wire          tg4_0_axi_rready;                                 // tg4_0:rready -> hbm_0_example_design:axi_4_0_rready
	wire    [7:0] tg4_0_axi_awlen;                                  // tg4_0:awlen -> hbm_0_example_design:axi_4_0_awlen
	wire    [3:0] tg4_0_axi_awqos;                                  // tg4_0:awqos -> hbm_0_example_design:axi_4_0_awqos
	wire          tg4_0_axi_wvalid;                                 // tg4_0:wvalid -> hbm_0_example_design:axi_4_0_wvalid
	wire   [29:0] tg4_0_axi_araddr;                                 // tg4_0:araddr -> hbm_0_example_design:axi_4_0_araddr
	wire    [2:0] tg4_0_axi_arprot;                                 // tg4_0:arprot -> hbm_0_example_design:axi_4_0_arprot
	wire    [2:0] tg4_0_axi_awprot;                                 // tg4_0:awprot -> hbm_0_example_design:axi_4_0_awprot
	wire  [255:0] tg4_0_axi_wdata;                                  // tg4_0:wdata -> hbm_0_example_design:axi_4_0_wdata
	wire          tg4_0_axi_arvalid;                                // tg4_0:arvalid -> hbm_0_example_design:axi_4_0_arvalid
	wire    [6:0] tg4_0_axi_arid;                                   // tg4_0:arid -> hbm_0_example_design:axi_4_0_arid
	wire   [29:0] tg4_0_axi_awaddr;                                 // tg4_0:awaddr -> hbm_0_example_design:axi_4_0_awaddr
	wire    [1:0] tg4_0_axi_bresp;                                  // hbm_0_example_design:axi_4_0_bresp -> tg4_0:bresp
	wire          tg4_0_axi_arready;                                // hbm_0_example_design:axi_4_0_arready -> tg4_0:arready
	wire  [255:0] tg4_0_axi_rdata;                                  // hbm_0_example_design:axi_4_0_rdata -> tg4_0:rdata
	wire          tg4_0_axi_awready;                                // hbm_0_example_design:axi_4_0_awready -> tg4_0:awready
	wire    [1:0] tg4_0_axi_arburst;                                // tg4_0:arburst -> hbm_0_example_design:axi_4_0_arburst
	wire    [2:0] tg4_0_axi_arsize;                                 // tg4_0:arsize -> hbm_0_example_design:axi_4_0_arsize
	wire          tg4_0_axi_bready;                                 // tg4_0:bready -> hbm_0_example_design:axi_4_0_bready
	wire          tg4_0_axi_rlast;                                  // hbm_0_example_design:axi_4_0_rlast -> tg4_0:rlast
	wire          tg4_0_axi_wlast;                                  // tg4_0:wlast -> hbm_0_example_design:axi_4_0_wlast
	wire    [1:0] tg4_0_axi_rresp;                                  // hbm_0_example_design:axi_4_0_rresp -> tg4_0:rresp
	wire    [6:0] tg4_0_axi_awid;                                   // tg4_0:awid -> hbm_0_example_design:axi_4_0_awid
	wire    [6:0] tg4_0_axi_bid;                                    // hbm_0_example_design:axi_4_0_bid -> tg4_0:bid
	wire          tg4_0_axi_bvalid;                                 // hbm_0_example_design:axi_4_0_bvalid -> tg4_0:bvalid
	wire    [2:0] tg4_0_axi_awsize;                                 // tg4_0:awsize -> hbm_0_example_design:axi_4_0_awsize
	wire          tg4_0_axi_awvalid;                                // tg4_0:awvalid -> hbm_0_example_design:axi_4_0_awvalid
	wire    [0:0] tg4_0_axi_aruser;                                 // tg4_0:aruser_ap -> hbm_0_example_design:axi_4_0_aruser
	wire          tg4_0_axi_rvalid;                                 // hbm_0_example_design:axi_4_0_rvalid -> tg4_0:rvalid
	wire    [1:0] tg4_1_axi_awburst;                                // tg4_1:awburst -> hbm_0_example_design:axi_4_1_awburst
	wire    [0:0] tg4_1_axi_awuser;                                 // tg4_1:awuser_ap -> hbm_0_example_design:axi_4_1_awuser
	wire    [7:0] tg4_1_axi_arlen;                                  // tg4_1:arlen -> hbm_0_example_design:axi_4_1_arlen
	wire    [3:0] tg4_1_axi_arqos;                                  // tg4_1:arqos -> hbm_0_example_design:axi_4_1_arqos
	wire   [31:0] tg4_1_axi_wstrb;                                  // tg4_1:wstrb -> hbm_0_example_design:axi_4_1_wstrb
	wire          tg4_1_axi_wready;                                 // hbm_0_example_design:axi_4_1_wready -> tg4_1:wready
	wire    [6:0] tg4_1_axi_rid;                                    // hbm_0_example_design:axi_4_1_rid -> tg4_1:rid
	wire          tg4_1_axi_rready;                                 // tg4_1:rready -> hbm_0_example_design:axi_4_1_rready
	wire    [7:0] tg4_1_axi_awlen;                                  // tg4_1:awlen -> hbm_0_example_design:axi_4_1_awlen
	wire    [3:0] tg4_1_axi_awqos;                                  // tg4_1:awqos -> hbm_0_example_design:axi_4_1_awqos
	wire          tg4_1_axi_wvalid;                                 // tg4_1:wvalid -> hbm_0_example_design:axi_4_1_wvalid
	wire   [29:0] tg4_1_axi_araddr;                                 // tg4_1:araddr -> hbm_0_example_design:axi_4_1_araddr
	wire    [2:0] tg4_1_axi_arprot;                                 // tg4_1:arprot -> hbm_0_example_design:axi_4_1_arprot
	wire    [2:0] tg4_1_axi_awprot;                                 // tg4_1:awprot -> hbm_0_example_design:axi_4_1_awprot
	wire  [255:0] tg4_1_axi_wdata;                                  // tg4_1:wdata -> hbm_0_example_design:axi_4_1_wdata
	wire          tg4_1_axi_arvalid;                                // tg4_1:arvalid -> hbm_0_example_design:axi_4_1_arvalid
	wire    [6:0] tg4_1_axi_arid;                                   // tg4_1:arid -> hbm_0_example_design:axi_4_1_arid
	wire   [29:0] tg4_1_axi_awaddr;                                 // tg4_1:awaddr -> hbm_0_example_design:axi_4_1_awaddr
	wire    [1:0] tg4_1_axi_bresp;                                  // hbm_0_example_design:axi_4_1_bresp -> tg4_1:bresp
	wire          tg4_1_axi_arready;                                // hbm_0_example_design:axi_4_1_arready -> tg4_1:arready
	wire  [255:0] tg4_1_axi_rdata;                                  // hbm_0_example_design:axi_4_1_rdata -> tg4_1:rdata
	wire          tg4_1_axi_awready;                                // hbm_0_example_design:axi_4_1_awready -> tg4_1:awready
	wire    [1:0] tg4_1_axi_arburst;                                // tg4_1:arburst -> hbm_0_example_design:axi_4_1_arburst
	wire    [2:0] tg4_1_axi_arsize;                                 // tg4_1:arsize -> hbm_0_example_design:axi_4_1_arsize
	wire          tg4_1_axi_bready;                                 // tg4_1:bready -> hbm_0_example_design:axi_4_1_bready
	wire          tg4_1_axi_rlast;                                  // hbm_0_example_design:axi_4_1_rlast -> tg4_1:rlast
	wire          tg4_1_axi_wlast;                                  // tg4_1:wlast -> hbm_0_example_design:axi_4_1_wlast
	wire    [1:0] tg4_1_axi_rresp;                                  // hbm_0_example_design:axi_4_1_rresp -> tg4_1:rresp
	wire    [6:0] tg4_1_axi_awid;                                   // tg4_1:awid -> hbm_0_example_design:axi_4_1_awid
	wire    [6:0] tg4_1_axi_bid;                                    // hbm_0_example_design:axi_4_1_bid -> tg4_1:bid
	wire          tg4_1_axi_bvalid;                                 // hbm_0_example_design:axi_4_1_bvalid -> tg4_1:bvalid
	wire    [2:0] tg4_1_axi_awsize;                                 // tg4_1:awsize -> hbm_0_example_design:axi_4_1_awsize
	wire          tg4_1_axi_awvalid;                                // tg4_1:awvalid -> hbm_0_example_design:axi_4_1_awvalid
	wire    [0:0] tg4_1_axi_aruser;                                 // tg4_1:aruser_ap -> hbm_0_example_design:axi_4_1_aruser
	wire          tg4_1_axi_rvalid;                                 // hbm_0_example_design:axi_4_1_rvalid -> tg4_1:rvalid
	wire    [1:0] tg5_0_axi_awburst;                                // tg5_0:awburst -> hbm_0_example_design:axi_5_0_awburst
	wire    [0:0] tg5_0_axi_awuser;                                 // tg5_0:awuser_ap -> hbm_0_example_design:axi_5_0_awuser
	wire    [7:0] tg5_0_axi_arlen;                                  // tg5_0:arlen -> hbm_0_example_design:axi_5_0_arlen
	wire    [3:0] tg5_0_axi_arqos;                                  // tg5_0:arqos -> hbm_0_example_design:axi_5_0_arqos
	wire   [31:0] tg5_0_axi_wstrb;                                  // tg5_0:wstrb -> hbm_0_example_design:axi_5_0_wstrb
	wire          tg5_0_axi_wready;                                 // hbm_0_example_design:axi_5_0_wready -> tg5_0:wready
	wire    [6:0] tg5_0_axi_rid;                                    // hbm_0_example_design:axi_5_0_rid -> tg5_0:rid
	wire          tg5_0_axi_rready;                                 // tg5_0:rready -> hbm_0_example_design:axi_5_0_rready
	wire    [7:0] tg5_0_axi_awlen;                                  // tg5_0:awlen -> hbm_0_example_design:axi_5_0_awlen
	wire    [3:0] tg5_0_axi_awqos;                                  // tg5_0:awqos -> hbm_0_example_design:axi_5_0_awqos
	wire          tg5_0_axi_wvalid;                                 // tg5_0:wvalid -> hbm_0_example_design:axi_5_0_wvalid
	wire   [29:0] tg5_0_axi_araddr;                                 // tg5_0:araddr -> hbm_0_example_design:axi_5_0_araddr
	wire    [2:0] tg5_0_axi_arprot;                                 // tg5_0:arprot -> hbm_0_example_design:axi_5_0_arprot
	wire    [2:0] tg5_0_axi_awprot;                                 // tg5_0:awprot -> hbm_0_example_design:axi_5_0_awprot
	wire  [255:0] tg5_0_axi_wdata;                                  // tg5_0:wdata -> hbm_0_example_design:axi_5_0_wdata
	wire          tg5_0_axi_arvalid;                                // tg5_0:arvalid -> hbm_0_example_design:axi_5_0_arvalid
	wire    [6:0] tg5_0_axi_arid;                                   // tg5_0:arid -> hbm_0_example_design:axi_5_0_arid
	wire   [29:0] tg5_0_axi_awaddr;                                 // tg5_0:awaddr -> hbm_0_example_design:axi_5_0_awaddr
	wire    [1:0] tg5_0_axi_bresp;                                  // hbm_0_example_design:axi_5_0_bresp -> tg5_0:bresp
	wire          tg5_0_axi_arready;                                // hbm_0_example_design:axi_5_0_arready -> tg5_0:arready
	wire  [255:0] tg5_0_axi_rdata;                                  // hbm_0_example_design:axi_5_0_rdata -> tg5_0:rdata
	wire          tg5_0_axi_awready;                                // hbm_0_example_design:axi_5_0_awready -> tg5_0:awready
	wire    [1:0] tg5_0_axi_arburst;                                // tg5_0:arburst -> hbm_0_example_design:axi_5_0_arburst
	wire    [2:0] tg5_0_axi_arsize;                                 // tg5_0:arsize -> hbm_0_example_design:axi_5_0_arsize
	wire          tg5_0_axi_bready;                                 // tg5_0:bready -> hbm_0_example_design:axi_5_0_bready
	wire          tg5_0_axi_rlast;                                  // hbm_0_example_design:axi_5_0_rlast -> tg5_0:rlast
	wire          tg5_0_axi_wlast;                                  // tg5_0:wlast -> hbm_0_example_design:axi_5_0_wlast
	wire    [1:0] tg5_0_axi_rresp;                                  // hbm_0_example_design:axi_5_0_rresp -> tg5_0:rresp
	wire    [6:0] tg5_0_axi_awid;                                   // tg5_0:awid -> hbm_0_example_design:axi_5_0_awid
	wire    [6:0] tg5_0_axi_bid;                                    // hbm_0_example_design:axi_5_0_bid -> tg5_0:bid
	wire          tg5_0_axi_bvalid;                                 // hbm_0_example_design:axi_5_0_bvalid -> tg5_0:bvalid
	wire    [2:0] tg5_0_axi_awsize;                                 // tg5_0:awsize -> hbm_0_example_design:axi_5_0_awsize
	wire          tg5_0_axi_awvalid;                                // tg5_0:awvalid -> hbm_0_example_design:axi_5_0_awvalid
	wire    [0:0] tg5_0_axi_aruser;                                 // tg5_0:aruser_ap -> hbm_0_example_design:axi_5_0_aruser
	wire          tg5_0_axi_rvalid;                                 // hbm_0_example_design:axi_5_0_rvalid -> tg5_0:rvalid
	wire    [1:0] tg5_1_axi_awburst;                                // tg5_1:awburst -> hbm_0_example_design:axi_5_1_awburst
	wire    [0:0] tg5_1_axi_awuser;                                 // tg5_1:awuser_ap -> hbm_0_example_design:axi_5_1_awuser
	wire    [7:0] tg5_1_axi_arlen;                                  // tg5_1:arlen -> hbm_0_example_design:axi_5_1_arlen
	wire    [3:0] tg5_1_axi_arqos;                                  // tg5_1:arqos -> hbm_0_example_design:axi_5_1_arqos
	wire   [31:0] tg5_1_axi_wstrb;                                  // tg5_1:wstrb -> hbm_0_example_design:axi_5_1_wstrb
	wire          tg5_1_axi_wready;                                 // hbm_0_example_design:axi_5_1_wready -> tg5_1:wready
	wire    [6:0] tg5_1_axi_rid;                                    // hbm_0_example_design:axi_5_1_rid -> tg5_1:rid
	wire          tg5_1_axi_rready;                                 // tg5_1:rready -> hbm_0_example_design:axi_5_1_rready
	wire    [7:0] tg5_1_axi_awlen;                                  // tg5_1:awlen -> hbm_0_example_design:axi_5_1_awlen
	wire    [3:0] tg5_1_axi_awqos;                                  // tg5_1:awqos -> hbm_0_example_design:axi_5_1_awqos
	wire          tg5_1_axi_wvalid;                                 // tg5_1:wvalid -> hbm_0_example_design:axi_5_1_wvalid
	wire   [29:0] tg5_1_axi_araddr;                                 // tg5_1:araddr -> hbm_0_example_design:axi_5_1_araddr
	wire    [2:0] tg5_1_axi_arprot;                                 // tg5_1:arprot -> hbm_0_example_design:axi_5_1_arprot
	wire    [2:0] tg5_1_axi_awprot;                                 // tg5_1:awprot -> hbm_0_example_design:axi_5_1_awprot
	wire  [255:0] tg5_1_axi_wdata;                                  // tg5_1:wdata -> hbm_0_example_design:axi_5_1_wdata
	wire          tg5_1_axi_arvalid;                                // tg5_1:arvalid -> hbm_0_example_design:axi_5_1_arvalid
	wire    [6:0] tg5_1_axi_arid;                                   // tg5_1:arid -> hbm_0_example_design:axi_5_1_arid
	wire   [29:0] tg5_1_axi_awaddr;                                 // tg5_1:awaddr -> hbm_0_example_design:axi_5_1_awaddr
	wire    [1:0] tg5_1_axi_bresp;                                  // hbm_0_example_design:axi_5_1_bresp -> tg5_1:bresp
	wire          tg5_1_axi_arready;                                // hbm_0_example_design:axi_5_1_arready -> tg5_1:arready
	wire  [255:0] tg5_1_axi_rdata;                                  // hbm_0_example_design:axi_5_1_rdata -> tg5_1:rdata
	wire          tg5_1_axi_awready;                                // hbm_0_example_design:axi_5_1_awready -> tg5_1:awready
	wire    [1:0] tg5_1_axi_arburst;                                // tg5_1:arburst -> hbm_0_example_design:axi_5_1_arburst
	wire    [2:0] tg5_1_axi_arsize;                                 // tg5_1:arsize -> hbm_0_example_design:axi_5_1_arsize
	wire          tg5_1_axi_bready;                                 // tg5_1:bready -> hbm_0_example_design:axi_5_1_bready
	wire          tg5_1_axi_rlast;                                  // hbm_0_example_design:axi_5_1_rlast -> tg5_1:rlast
	wire          tg5_1_axi_wlast;                                  // tg5_1:wlast -> hbm_0_example_design:axi_5_1_wlast
	wire    [1:0] tg5_1_axi_rresp;                                  // hbm_0_example_design:axi_5_1_rresp -> tg5_1:rresp
	wire    [6:0] tg5_1_axi_awid;                                   // tg5_1:awid -> hbm_0_example_design:axi_5_1_awid
	wire    [6:0] tg5_1_axi_bid;                                    // hbm_0_example_design:axi_5_1_bid -> tg5_1:bid
	wire          tg5_1_axi_bvalid;                                 // hbm_0_example_design:axi_5_1_bvalid -> tg5_1:bvalid
	wire    [2:0] tg5_1_axi_awsize;                                 // tg5_1:awsize -> hbm_0_example_design:axi_5_1_awsize
	wire          tg5_1_axi_awvalid;                                // tg5_1:awvalid -> hbm_0_example_design:axi_5_1_awvalid
	wire    [0:0] tg5_1_axi_aruser;                                 // tg5_1:aruser_ap -> hbm_0_example_design:axi_5_1_aruser
	wire          tg5_1_axi_rvalid;                                 // hbm_0_example_design:axi_5_1_rvalid -> tg5_1:rvalid
	wire    [1:0] tg6_0_axi_awburst;                                // tg6_0:awburst -> hbm_0_example_design:axi_6_0_awburst
	wire    [0:0] tg6_0_axi_awuser;                                 // tg6_0:awuser_ap -> hbm_0_example_design:axi_6_0_awuser
	wire    [7:0] tg6_0_axi_arlen;                                  // tg6_0:arlen -> hbm_0_example_design:axi_6_0_arlen
	wire    [3:0] tg6_0_axi_arqos;                                  // tg6_0:arqos -> hbm_0_example_design:axi_6_0_arqos
	wire   [31:0] tg6_0_axi_wstrb;                                  // tg6_0:wstrb -> hbm_0_example_design:axi_6_0_wstrb
	wire          tg6_0_axi_wready;                                 // hbm_0_example_design:axi_6_0_wready -> tg6_0:wready
	wire    [6:0] tg6_0_axi_rid;                                    // hbm_0_example_design:axi_6_0_rid -> tg6_0:rid
	wire          tg6_0_axi_rready;                                 // tg6_0:rready -> hbm_0_example_design:axi_6_0_rready
	wire    [7:0] tg6_0_axi_awlen;                                  // tg6_0:awlen -> hbm_0_example_design:axi_6_0_awlen
	wire    [3:0] tg6_0_axi_awqos;                                  // tg6_0:awqos -> hbm_0_example_design:axi_6_0_awqos
	wire          tg6_0_axi_wvalid;                                 // tg6_0:wvalid -> hbm_0_example_design:axi_6_0_wvalid
	wire   [29:0] tg6_0_axi_araddr;                                 // tg6_0:araddr -> hbm_0_example_design:axi_6_0_araddr
	wire    [2:0] tg6_0_axi_arprot;                                 // tg6_0:arprot -> hbm_0_example_design:axi_6_0_arprot
	wire    [2:0] tg6_0_axi_awprot;                                 // tg6_0:awprot -> hbm_0_example_design:axi_6_0_awprot
	wire  [255:0] tg6_0_axi_wdata;                                  // tg6_0:wdata -> hbm_0_example_design:axi_6_0_wdata
	wire          tg6_0_axi_arvalid;                                // tg6_0:arvalid -> hbm_0_example_design:axi_6_0_arvalid
	wire    [6:0] tg6_0_axi_arid;                                   // tg6_0:arid -> hbm_0_example_design:axi_6_0_arid
	wire   [29:0] tg6_0_axi_awaddr;                                 // tg6_0:awaddr -> hbm_0_example_design:axi_6_0_awaddr
	wire    [1:0] tg6_0_axi_bresp;                                  // hbm_0_example_design:axi_6_0_bresp -> tg6_0:bresp
	wire          tg6_0_axi_arready;                                // hbm_0_example_design:axi_6_0_arready -> tg6_0:arready
	wire  [255:0] tg6_0_axi_rdata;                                  // hbm_0_example_design:axi_6_0_rdata -> tg6_0:rdata
	wire          tg6_0_axi_awready;                                // hbm_0_example_design:axi_6_0_awready -> tg6_0:awready
	wire    [1:0] tg6_0_axi_arburst;                                // tg6_0:arburst -> hbm_0_example_design:axi_6_0_arburst
	wire    [2:0] tg6_0_axi_arsize;                                 // tg6_0:arsize -> hbm_0_example_design:axi_6_0_arsize
	wire          tg6_0_axi_bready;                                 // tg6_0:bready -> hbm_0_example_design:axi_6_0_bready
	wire          tg6_0_axi_rlast;                                  // hbm_0_example_design:axi_6_0_rlast -> tg6_0:rlast
	wire          tg6_0_axi_wlast;                                  // tg6_0:wlast -> hbm_0_example_design:axi_6_0_wlast
	wire    [1:0] tg6_0_axi_rresp;                                  // hbm_0_example_design:axi_6_0_rresp -> tg6_0:rresp
	wire    [6:0] tg6_0_axi_awid;                                   // tg6_0:awid -> hbm_0_example_design:axi_6_0_awid
	wire    [6:0] tg6_0_axi_bid;                                    // hbm_0_example_design:axi_6_0_bid -> tg6_0:bid
	wire          tg6_0_axi_bvalid;                                 // hbm_0_example_design:axi_6_0_bvalid -> tg6_0:bvalid
	wire    [2:0] tg6_0_axi_awsize;                                 // tg6_0:awsize -> hbm_0_example_design:axi_6_0_awsize
	wire          tg6_0_axi_awvalid;                                // tg6_0:awvalid -> hbm_0_example_design:axi_6_0_awvalid
	wire    [0:0] tg6_0_axi_aruser;                                 // tg6_0:aruser_ap -> hbm_0_example_design:axi_6_0_aruser
	wire          tg6_0_axi_rvalid;                                 // hbm_0_example_design:axi_6_0_rvalid -> tg6_0:rvalid
	wire    [1:0] tg6_1_axi_awburst;                                // tg6_1:awburst -> hbm_0_example_design:axi_6_1_awburst
	wire    [0:0] tg6_1_axi_awuser;                                 // tg6_1:awuser_ap -> hbm_0_example_design:axi_6_1_awuser
	wire    [7:0] tg6_1_axi_arlen;                                  // tg6_1:arlen -> hbm_0_example_design:axi_6_1_arlen
	wire    [3:0] tg6_1_axi_arqos;                                  // tg6_1:arqos -> hbm_0_example_design:axi_6_1_arqos
	wire   [31:0] tg6_1_axi_wstrb;                                  // tg6_1:wstrb -> hbm_0_example_design:axi_6_1_wstrb
	wire          tg6_1_axi_wready;                                 // hbm_0_example_design:axi_6_1_wready -> tg6_1:wready
	wire    [6:0] tg6_1_axi_rid;                                    // hbm_0_example_design:axi_6_1_rid -> tg6_1:rid
	wire          tg6_1_axi_rready;                                 // tg6_1:rready -> hbm_0_example_design:axi_6_1_rready
	wire    [7:0] tg6_1_axi_awlen;                                  // tg6_1:awlen -> hbm_0_example_design:axi_6_1_awlen
	wire    [3:0] tg6_1_axi_awqos;                                  // tg6_1:awqos -> hbm_0_example_design:axi_6_1_awqos
	wire          tg6_1_axi_wvalid;                                 // tg6_1:wvalid -> hbm_0_example_design:axi_6_1_wvalid
	wire   [29:0] tg6_1_axi_araddr;                                 // tg6_1:araddr -> hbm_0_example_design:axi_6_1_araddr
	wire    [2:0] tg6_1_axi_arprot;                                 // tg6_1:arprot -> hbm_0_example_design:axi_6_1_arprot
	wire    [2:0] tg6_1_axi_awprot;                                 // tg6_1:awprot -> hbm_0_example_design:axi_6_1_awprot
	wire  [255:0] tg6_1_axi_wdata;                                  // tg6_1:wdata -> hbm_0_example_design:axi_6_1_wdata
	wire          tg6_1_axi_arvalid;                                // tg6_1:arvalid -> hbm_0_example_design:axi_6_1_arvalid
	wire    [6:0] tg6_1_axi_arid;                                   // tg6_1:arid -> hbm_0_example_design:axi_6_1_arid
	wire   [29:0] tg6_1_axi_awaddr;                                 // tg6_1:awaddr -> hbm_0_example_design:axi_6_1_awaddr
	wire    [1:0] tg6_1_axi_bresp;                                  // hbm_0_example_design:axi_6_1_bresp -> tg6_1:bresp
	wire          tg6_1_axi_arready;                                // hbm_0_example_design:axi_6_1_arready -> tg6_1:arready
	wire  [255:0] tg6_1_axi_rdata;                                  // hbm_0_example_design:axi_6_1_rdata -> tg6_1:rdata
	wire          tg6_1_axi_awready;                                // hbm_0_example_design:axi_6_1_awready -> tg6_1:awready
	wire    [1:0] tg6_1_axi_arburst;                                // tg6_1:arburst -> hbm_0_example_design:axi_6_1_arburst
	wire    [2:0] tg6_1_axi_arsize;                                 // tg6_1:arsize -> hbm_0_example_design:axi_6_1_arsize
	wire          tg6_1_axi_bready;                                 // tg6_1:bready -> hbm_0_example_design:axi_6_1_bready
	wire          tg6_1_axi_rlast;                                  // hbm_0_example_design:axi_6_1_rlast -> tg6_1:rlast
	wire          tg6_1_axi_wlast;                                  // tg6_1:wlast -> hbm_0_example_design:axi_6_1_wlast
	wire    [1:0] tg6_1_axi_rresp;                                  // hbm_0_example_design:axi_6_1_rresp -> tg6_1:rresp
	wire    [6:0] tg6_1_axi_awid;                                   // tg6_1:awid -> hbm_0_example_design:axi_6_1_awid
	wire    [6:0] tg6_1_axi_bid;                                    // hbm_0_example_design:axi_6_1_bid -> tg6_1:bid
	wire          tg6_1_axi_bvalid;                                 // hbm_0_example_design:axi_6_1_bvalid -> tg6_1:bvalid
	wire    [2:0] tg6_1_axi_awsize;                                 // tg6_1:awsize -> hbm_0_example_design:axi_6_1_awsize
	wire          tg6_1_axi_awvalid;                                // tg6_1:awvalid -> hbm_0_example_design:axi_6_1_awvalid
	wire    [0:0] tg6_1_axi_aruser;                                 // tg6_1:aruser_ap -> hbm_0_example_design:axi_6_1_aruser
	wire          tg6_1_axi_rvalid;                                 // hbm_0_example_design:axi_6_1_rvalid -> tg6_1:rvalid
	wire    [1:0] tg7_0_axi_awburst;                                // tg7_0:awburst -> hbm_0_example_design:axi_7_0_awburst
	wire    [0:0] tg7_0_axi_awuser;                                 // tg7_0:awuser_ap -> hbm_0_example_design:axi_7_0_awuser
	wire    [7:0] tg7_0_axi_arlen;                                  // tg7_0:arlen -> hbm_0_example_design:axi_7_0_arlen
	wire    [3:0] tg7_0_axi_arqos;                                  // tg7_0:arqos -> hbm_0_example_design:axi_7_0_arqos
	wire   [31:0] tg7_0_axi_wstrb;                                  // tg7_0:wstrb -> hbm_0_example_design:axi_7_0_wstrb
	wire          tg7_0_axi_wready;                                 // hbm_0_example_design:axi_7_0_wready -> tg7_0:wready
	wire    [6:0] tg7_0_axi_rid;                                    // hbm_0_example_design:axi_7_0_rid -> tg7_0:rid
	wire          tg7_0_axi_rready;                                 // tg7_0:rready -> hbm_0_example_design:axi_7_0_rready
	wire    [7:0] tg7_0_axi_awlen;                                  // tg7_0:awlen -> hbm_0_example_design:axi_7_0_awlen
	wire    [3:0] tg7_0_axi_awqos;                                  // tg7_0:awqos -> hbm_0_example_design:axi_7_0_awqos
	wire          tg7_0_axi_wvalid;                                 // tg7_0:wvalid -> hbm_0_example_design:axi_7_0_wvalid
	wire   [29:0] tg7_0_axi_araddr;                                 // tg7_0:araddr -> hbm_0_example_design:axi_7_0_araddr
	wire    [2:0] tg7_0_axi_arprot;                                 // tg7_0:arprot -> hbm_0_example_design:axi_7_0_arprot
	wire    [2:0] tg7_0_axi_awprot;                                 // tg7_0:awprot -> hbm_0_example_design:axi_7_0_awprot
	wire  [255:0] tg7_0_axi_wdata;                                  // tg7_0:wdata -> hbm_0_example_design:axi_7_0_wdata
	wire          tg7_0_axi_arvalid;                                // tg7_0:arvalid -> hbm_0_example_design:axi_7_0_arvalid
	wire    [6:0] tg7_0_axi_arid;                                   // tg7_0:arid -> hbm_0_example_design:axi_7_0_arid
	wire   [29:0] tg7_0_axi_awaddr;                                 // tg7_0:awaddr -> hbm_0_example_design:axi_7_0_awaddr
	wire    [1:0] tg7_0_axi_bresp;                                  // hbm_0_example_design:axi_7_0_bresp -> tg7_0:bresp
	wire          tg7_0_axi_arready;                                // hbm_0_example_design:axi_7_0_arready -> tg7_0:arready
	wire  [255:0] tg7_0_axi_rdata;                                  // hbm_0_example_design:axi_7_0_rdata -> tg7_0:rdata
	wire          tg7_0_axi_awready;                                // hbm_0_example_design:axi_7_0_awready -> tg7_0:awready
	wire    [1:0] tg7_0_axi_arburst;                                // tg7_0:arburst -> hbm_0_example_design:axi_7_0_arburst
	wire    [2:0] tg7_0_axi_arsize;                                 // tg7_0:arsize -> hbm_0_example_design:axi_7_0_arsize
	wire          tg7_0_axi_bready;                                 // tg7_0:bready -> hbm_0_example_design:axi_7_0_bready
	wire          tg7_0_axi_rlast;                                  // hbm_0_example_design:axi_7_0_rlast -> tg7_0:rlast
	wire          tg7_0_axi_wlast;                                  // tg7_0:wlast -> hbm_0_example_design:axi_7_0_wlast
	wire    [1:0] tg7_0_axi_rresp;                                  // hbm_0_example_design:axi_7_0_rresp -> tg7_0:rresp
	wire    [6:0] tg7_0_axi_awid;                                   // tg7_0:awid -> hbm_0_example_design:axi_7_0_awid
	wire    [6:0] tg7_0_axi_bid;                                    // hbm_0_example_design:axi_7_0_bid -> tg7_0:bid
	wire          tg7_0_axi_bvalid;                                 // hbm_0_example_design:axi_7_0_bvalid -> tg7_0:bvalid
	wire    [2:0] tg7_0_axi_awsize;                                 // tg7_0:awsize -> hbm_0_example_design:axi_7_0_awsize
	wire          tg7_0_axi_awvalid;                                // tg7_0:awvalid -> hbm_0_example_design:axi_7_0_awvalid
	wire    [0:0] tg7_0_axi_aruser;                                 // tg7_0:aruser_ap -> hbm_0_example_design:axi_7_0_aruser
	wire          tg7_0_axi_rvalid;                                 // hbm_0_example_design:axi_7_0_rvalid -> tg7_0:rvalid
	wire    [1:0] tg7_1_axi_awburst;                                // tg7_1:awburst -> hbm_0_example_design:axi_7_1_awburst
	wire    [0:0] tg7_1_axi_awuser;                                 // tg7_1:awuser_ap -> hbm_0_example_design:axi_7_1_awuser
	wire    [7:0] tg7_1_axi_arlen;                                  // tg7_1:arlen -> hbm_0_example_design:axi_7_1_arlen
	wire    [3:0] tg7_1_axi_arqos;                                  // tg7_1:arqos -> hbm_0_example_design:axi_7_1_arqos
	wire   [31:0] tg7_1_axi_wstrb;                                  // tg7_1:wstrb -> hbm_0_example_design:axi_7_1_wstrb
	wire          tg7_1_axi_wready;                                 // hbm_0_example_design:axi_7_1_wready -> tg7_1:wready
	wire    [6:0] tg7_1_axi_rid;                                    // hbm_0_example_design:axi_7_1_rid -> tg7_1:rid
	wire          tg7_1_axi_rready;                                 // tg7_1:rready -> hbm_0_example_design:axi_7_1_rready
	wire    [7:0] tg7_1_axi_awlen;                                  // tg7_1:awlen -> hbm_0_example_design:axi_7_1_awlen
	wire    [3:0] tg7_1_axi_awqos;                                  // tg7_1:awqos -> hbm_0_example_design:axi_7_1_awqos
	wire          tg7_1_axi_wvalid;                                 // tg7_1:wvalid -> hbm_0_example_design:axi_7_1_wvalid
	wire   [29:0] tg7_1_axi_araddr;                                 // tg7_1:araddr -> hbm_0_example_design:axi_7_1_araddr
	wire    [2:0] tg7_1_axi_arprot;                                 // tg7_1:arprot -> hbm_0_example_design:axi_7_1_arprot
	wire    [2:0] tg7_1_axi_awprot;                                 // tg7_1:awprot -> hbm_0_example_design:axi_7_1_awprot
	wire  [255:0] tg7_1_axi_wdata;                                  // tg7_1:wdata -> hbm_0_example_design:axi_7_1_wdata
	wire          tg7_1_axi_arvalid;                                // tg7_1:arvalid -> hbm_0_example_design:axi_7_1_arvalid
	wire    [6:0] tg7_1_axi_arid;                                   // tg7_1:arid -> hbm_0_example_design:axi_7_1_arid
	wire   [29:0] tg7_1_axi_awaddr;                                 // tg7_1:awaddr -> hbm_0_example_design:axi_7_1_awaddr
	wire    [1:0] tg7_1_axi_bresp;                                  // hbm_0_example_design:axi_7_1_bresp -> tg7_1:bresp
	wire          tg7_1_axi_arready;                                // hbm_0_example_design:axi_7_1_arready -> tg7_1:arready
	wire  [255:0] tg7_1_axi_rdata;                                  // hbm_0_example_design:axi_7_1_rdata -> tg7_1:rdata
	wire          tg7_1_axi_awready;                                // hbm_0_example_design:axi_7_1_awready -> tg7_1:awready
	wire    [1:0] tg7_1_axi_arburst;                                // tg7_1:arburst -> hbm_0_example_design:axi_7_1_arburst
	wire    [2:0] tg7_1_axi_arsize;                                 // tg7_1:arsize -> hbm_0_example_design:axi_7_1_arsize
	wire          tg7_1_axi_bready;                                 // tg7_1:bready -> hbm_0_example_design:axi_7_1_bready
	wire          tg7_1_axi_rlast;                                  // hbm_0_example_design:axi_7_1_rlast -> tg7_1:rlast
	wire          tg7_1_axi_wlast;                                  // tg7_1:wlast -> hbm_0_example_design:axi_7_1_wlast
	wire    [1:0] tg7_1_axi_rresp;                                  // hbm_0_example_design:axi_7_1_rresp -> tg7_1:rresp
	wire    [6:0] tg7_1_axi_awid;                                   // tg7_1:awid -> hbm_0_example_design:axi_7_1_awid
	wire    [6:0] tg7_1_axi_bid;                                    // hbm_0_example_design:axi_7_1_bid -> tg7_1:bid
	wire          tg7_1_axi_bvalid;                                 // hbm_0_example_design:axi_7_1_bvalid -> tg7_1:bvalid
	wire    [2:0] tg7_1_axi_awsize;                                 // tg7_1:awsize -> hbm_0_example_design:axi_7_1_awsize
	wire          tg7_1_axi_awvalid;                                // tg7_1:awvalid -> hbm_0_example_design:axi_7_1_awvalid
	wire    [0:0] tg7_1_axi_aruser;                                 // tg7_1:aruser_ap -> hbm_0_example_design:axi_7_1_aruser
	wire          tg7_1_axi_rvalid;                                 // hbm_0_example_design:axi_7_1_rvalid -> tg7_1:rvalid
	wire          core_clk_iopll_outclk0_clk;                       // core_clk_iopll:outclk_0 -> hbm_0_example_design:ext_core_clk
	wire          hbm_0_example_design_wmc_clk_0_clk;               // hbm_0_example_design:wmc_clk_0 -> [tg0_0:wmc_clk_in, tg0_1:wmc_clk_in, tg1_0:wmc_clk_in, tg1_1:wmc_clk_in]
	wire          hbm_0_example_design_wmc_clk_2_clk;               // hbm_0_example_design:wmc_clk_2 -> [tg2_0:wmc_clk_in, tg2_1:wmc_clk_in, tg3_0:wmc_clk_in, tg3_1:wmc_clk_in]
	wire          hbm_0_example_design_wmc_clk_4_clk;               // hbm_0_example_design:wmc_clk_4 -> [tg4_0:wmc_clk_in, tg4_1:wmc_clk_in, tg5_0:wmc_clk_in, tg5_1:wmc_clk_in]
	wire          hbm_0_example_design_wmc_clk_6_clk;               // hbm_0_example_design:wmc_clk_6 -> [tg6_0:wmc_clk_in, tg6_1:wmc_clk_in, tg7_0:wmc_clk_in, tg7_1:wmc_clk_in]
	wire    [1:0] tg0_0_apb_ur_pstrb;                               // tg0_0:ur_pstrb -> hbm_0_example_design:apb_0_ur_pstrb
	wire   [15:0] tg0_0_apb_ur_pwdata;                              // tg0_0:ur_pwdata -> hbm_0_example_design:apb_0_ur_pwdata
	wire          tg0_0_apb_ur_penable;                             // tg0_0:ur_penable -> hbm_0_example_design:apb_0_ur_penable
	wire   [15:0] tg0_0_apb_ur_paddr;                               // tg0_0:ur_paddr -> hbm_0_example_design:apb_0_ur_paddr
	wire          tg0_0_apb_ur_psel;                                // tg0_0:ur_psel -> hbm_0_example_design:apb_0_ur_psel
	wire          tg0_0_apb_ur_pwrite;                              // tg0_0:ur_pwrite -> hbm_0_example_design:apb_0_ur_pwrite
	wire          hbm_0_example_design_apb_0_ur_prready;            // hbm_0_example_design:apb_0_ur_prready -> tg0_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_0_ur_prdata;             // hbm_0_example_design:apb_0_ur_prdata -> tg0_0:ur_prdata
	wire    [1:0] tg1_0_apb_ur_pstrb;                               // tg1_0:ur_pstrb -> hbm_0_example_design:apb_1_ur_pstrb
	wire   [15:0] tg1_0_apb_ur_pwdata;                              // tg1_0:ur_pwdata -> hbm_0_example_design:apb_1_ur_pwdata
	wire          tg1_0_apb_ur_penable;                             // tg1_0:ur_penable -> hbm_0_example_design:apb_1_ur_penable
	wire   [15:0] tg1_0_apb_ur_paddr;                               // tg1_0:ur_paddr -> hbm_0_example_design:apb_1_ur_paddr
	wire          tg1_0_apb_ur_psel;                                // tg1_0:ur_psel -> hbm_0_example_design:apb_1_ur_psel
	wire          tg1_0_apb_ur_pwrite;                              // tg1_0:ur_pwrite -> hbm_0_example_design:apb_1_ur_pwrite
	wire          hbm_0_example_design_apb_1_ur_prready;            // hbm_0_example_design:apb_1_ur_prready -> tg1_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_1_ur_prdata;             // hbm_0_example_design:apb_1_ur_prdata -> tg1_0:ur_prdata
	wire    [1:0] tg2_0_apb_ur_pstrb;                               // tg2_0:ur_pstrb -> hbm_0_example_design:apb_2_ur_pstrb
	wire   [15:0] tg2_0_apb_ur_pwdata;                              // tg2_0:ur_pwdata -> hbm_0_example_design:apb_2_ur_pwdata
	wire          tg2_0_apb_ur_penable;                             // tg2_0:ur_penable -> hbm_0_example_design:apb_2_ur_penable
	wire   [15:0] tg2_0_apb_ur_paddr;                               // tg2_0:ur_paddr -> hbm_0_example_design:apb_2_ur_paddr
	wire          tg2_0_apb_ur_psel;                                // tg2_0:ur_psel -> hbm_0_example_design:apb_2_ur_psel
	wire          tg2_0_apb_ur_pwrite;                              // tg2_0:ur_pwrite -> hbm_0_example_design:apb_2_ur_pwrite
	wire          hbm_0_example_design_apb_2_ur_prready;            // hbm_0_example_design:apb_2_ur_prready -> tg2_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_2_ur_prdata;             // hbm_0_example_design:apb_2_ur_prdata -> tg2_0:ur_prdata
	wire    [1:0] tg3_0_apb_ur_pstrb;                               // tg3_0:ur_pstrb -> hbm_0_example_design:apb_3_ur_pstrb
	wire   [15:0] tg3_0_apb_ur_pwdata;                              // tg3_0:ur_pwdata -> hbm_0_example_design:apb_3_ur_pwdata
	wire          tg3_0_apb_ur_penable;                             // tg3_0:ur_penable -> hbm_0_example_design:apb_3_ur_penable
	wire   [15:0] tg3_0_apb_ur_paddr;                               // tg3_0:ur_paddr -> hbm_0_example_design:apb_3_ur_paddr
	wire          tg3_0_apb_ur_psel;                                // tg3_0:ur_psel -> hbm_0_example_design:apb_3_ur_psel
	wire          tg3_0_apb_ur_pwrite;                              // tg3_0:ur_pwrite -> hbm_0_example_design:apb_3_ur_pwrite
	wire          hbm_0_example_design_apb_3_ur_prready;            // hbm_0_example_design:apb_3_ur_prready -> tg3_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_3_ur_prdata;             // hbm_0_example_design:apb_3_ur_prdata -> tg3_0:ur_prdata
	wire    [1:0] tg4_0_apb_ur_pstrb;                               // tg4_0:ur_pstrb -> hbm_0_example_design:apb_4_ur_pstrb
	wire   [15:0] tg4_0_apb_ur_pwdata;                              // tg4_0:ur_pwdata -> hbm_0_example_design:apb_4_ur_pwdata
	wire          tg4_0_apb_ur_penable;                             // tg4_0:ur_penable -> hbm_0_example_design:apb_4_ur_penable
	wire   [15:0] tg4_0_apb_ur_paddr;                               // tg4_0:ur_paddr -> hbm_0_example_design:apb_4_ur_paddr
	wire          tg4_0_apb_ur_psel;                                // tg4_0:ur_psel -> hbm_0_example_design:apb_4_ur_psel
	wire          tg4_0_apb_ur_pwrite;                              // tg4_0:ur_pwrite -> hbm_0_example_design:apb_4_ur_pwrite
	wire          hbm_0_example_design_apb_4_ur_prready;            // hbm_0_example_design:apb_4_ur_prready -> tg4_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_4_ur_prdata;             // hbm_0_example_design:apb_4_ur_prdata -> tg4_0:ur_prdata
	wire    [1:0] tg5_0_apb_ur_pstrb;                               // tg5_0:ur_pstrb -> hbm_0_example_design:apb_5_ur_pstrb
	wire   [15:0] tg5_0_apb_ur_pwdata;                              // tg5_0:ur_pwdata -> hbm_0_example_design:apb_5_ur_pwdata
	wire          tg5_0_apb_ur_penable;                             // tg5_0:ur_penable -> hbm_0_example_design:apb_5_ur_penable
	wire   [15:0] tg5_0_apb_ur_paddr;                               // tg5_0:ur_paddr -> hbm_0_example_design:apb_5_ur_paddr
	wire          tg5_0_apb_ur_psel;                                // tg5_0:ur_psel -> hbm_0_example_design:apb_5_ur_psel
	wire          tg5_0_apb_ur_pwrite;                              // tg5_0:ur_pwrite -> hbm_0_example_design:apb_5_ur_pwrite
	wire          hbm_0_example_design_apb_5_ur_prready;            // hbm_0_example_design:apb_5_ur_prready -> tg5_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_5_ur_prdata;             // hbm_0_example_design:apb_5_ur_prdata -> tg5_0:ur_prdata
	wire    [1:0] tg6_0_apb_ur_pstrb;                               // tg6_0:ur_pstrb -> hbm_0_example_design:apb_6_ur_pstrb
	wire   [15:0] tg6_0_apb_ur_pwdata;                              // tg6_0:ur_pwdata -> hbm_0_example_design:apb_6_ur_pwdata
	wire          tg6_0_apb_ur_penable;                             // tg6_0:ur_penable -> hbm_0_example_design:apb_6_ur_penable
	wire   [15:0] tg6_0_apb_ur_paddr;                               // tg6_0:ur_paddr -> hbm_0_example_design:apb_6_ur_paddr
	wire          tg6_0_apb_ur_psel;                                // tg6_0:ur_psel -> hbm_0_example_design:apb_6_ur_psel
	wire          tg6_0_apb_ur_pwrite;                              // tg6_0:ur_pwrite -> hbm_0_example_design:apb_6_ur_pwrite
	wire          hbm_0_example_design_apb_6_ur_prready;            // hbm_0_example_design:apb_6_ur_prready -> tg6_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_6_ur_prdata;             // hbm_0_example_design:apb_6_ur_prdata -> tg6_0:ur_prdata
	wire    [1:0] tg7_0_apb_ur_pstrb;                               // tg7_0:ur_pstrb -> hbm_0_example_design:apb_7_ur_pstrb
	wire   [15:0] tg7_0_apb_ur_pwdata;                              // tg7_0:ur_pwdata -> hbm_0_example_design:apb_7_ur_pwdata
	wire          tg7_0_apb_ur_penable;                             // tg7_0:ur_penable -> hbm_0_example_design:apb_7_ur_penable
	wire   [15:0] tg7_0_apb_ur_paddr;                               // tg7_0:ur_paddr -> hbm_0_example_design:apb_7_ur_paddr
	wire          tg7_0_apb_ur_psel;                                // tg7_0:ur_psel -> hbm_0_example_design:apb_7_ur_psel
	wire          tg7_0_apb_ur_pwrite;                              // tg7_0:ur_pwrite -> hbm_0_example_design:apb_7_ur_pwrite
	wire          hbm_0_example_design_apb_7_ur_prready;            // hbm_0_example_design:apb_7_ur_prready -> tg7_0:ur_prready
	wire   [15:0] hbm_0_example_design_apb_7_ur_prdata;             // hbm_0_example_design:apb_7_ur_prdata -> tg7_0:ur_prdata
	wire          hbm_0_example_design_axi_extra_0_0_ruser_err_dbe; // hbm_0_example_design:axi_extra_0_0_ruser_err_dbe -> tg0_0:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_0_0_ruser_data;    // hbm_0_example_design:axi_extra_0_0_ruser_data -> tg0_0:ruser_data
	wire    [3:0] tg0_0_axi_extra_wuser_strb;                       // tg0_0:wuser_strb -> hbm_0_example_design:axi_extra_0_0_wuser_strb
	wire   [31:0] tg0_0_axi_extra_wuser_data;                       // tg0_0:wuser_data -> hbm_0_example_design:axi_extra_0_0_wuser_data
	wire          hbm_0_example_design_axi_extra_0_1_ruser_err_dbe; // hbm_0_example_design:axi_extra_0_1_ruser_err_dbe -> tg0_1:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_0_1_ruser_data;    // hbm_0_example_design:axi_extra_0_1_ruser_data -> tg0_1:ruser_data
	wire    [3:0] tg0_1_axi_extra_wuser_strb;                       // tg0_1:wuser_strb -> hbm_0_example_design:axi_extra_0_1_wuser_strb
	wire   [31:0] tg0_1_axi_extra_wuser_data;                       // tg0_1:wuser_data -> hbm_0_example_design:axi_extra_0_1_wuser_data
	wire          hbm_0_example_design_axi_extra_1_0_ruser_err_dbe; // hbm_0_example_design:axi_extra_1_0_ruser_err_dbe -> tg1_0:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_1_0_ruser_data;    // hbm_0_example_design:axi_extra_1_0_ruser_data -> tg1_0:ruser_data
	wire    [3:0] tg1_0_axi_extra_wuser_strb;                       // tg1_0:wuser_strb -> hbm_0_example_design:axi_extra_1_0_wuser_strb
	wire   [31:0] tg1_0_axi_extra_wuser_data;                       // tg1_0:wuser_data -> hbm_0_example_design:axi_extra_1_0_wuser_data
	wire          hbm_0_example_design_axi_extra_1_1_ruser_err_dbe; // hbm_0_example_design:axi_extra_1_1_ruser_err_dbe -> tg1_1:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_1_1_ruser_data;    // hbm_0_example_design:axi_extra_1_1_ruser_data -> tg1_1:ruser_data
	wire    [3:0] tg1_1_axi_extra_wuser_strb;                       // tg1_1:wuser_strb -> hbm_0_example_design:axi_extra_1_1_wuser_strb
	wire   [31:0] tg1_1_axi_extra_wuser_data;                       // tg1_1:wuser_data -> hbm_0_example_design:axi_extra_1_1_wuser_data
	wire          hbm_0_example_design_axi_extra_2_0_ruser_err_dbe; // hbm_0_example_design:axi_extra_2_0_ruser_err_dbe -> tg2_0:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_2_0_ruser_data;    // hbm_0_example_design:axi_extra_2_0_ruser_data -> tg2_0:ruser_data
	wire    [3:0] tg2_0_axi_extra_wuser_strb;                       // tg2_0:wuser_strb -> hbm_0_example_design:axi_extra_2_0_wuser_strb
	wire   [31:0] tg2_0_axi_extra_wuser_data;                       // tg2_0:wuser_data -> hbm_0_example_design:axi_extra_2_0_wuser_data
	wire          hbm_0_example_design_axi_extra_2_1_ruser_err_dbe; // hbm_0_example_design:axi_extra_2_1_ruser_err_dbe -> tg2_1:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_2_1_ruser_data;    // hbm_0_example_design:axi_extra_2_1_ruser_data -> tg2_1:ruser_data
	wire    [3:0] tg2_1_axi_extra_wuser_strb;                       // tg2_1:wuser_strb -> hbm_0_example_design:axi_extra_2_1_wuser_strb
	wire   [31:0] tg2_1_axi_extra_wuser_data;                       // tg2_1:wuser_data -> hbm_0_example_design:axi_extra_2_1_wuser_data
	wire          hbm_0_example_design_axi_extra_3_0_ruser_err_dbe; // hbm_0_example_design:axi_extra_3_0_ruser_err_dbe -> tg3_0:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_3_0_ruser_data;    // hbm_0_example_design:axi_extra_3_0_ruser_data -> tg3_0:ruser_data
	wire    [3:0] tg3_0_axi_extra_wuser_strb;                       // tg3_0:wuser_strb -> hbm_0_example_design:axi_extra_3_0_wuser_strb
	wire   [31:0] tg3_0_axi_extra_wuser_data;                       // tg3_0:wuser_data -> hbm_0_example_design:axi_extra_3_0_wuser_data
	wire          hbm_0_example_design_axi_extra_3_1_ruser_err_dbe; // hbm_0_example_design:axi_extra_3_1_ruser_err_dbe -> tg3_1:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_3_1_ruser_data;    // hbm_0_example_design:axi_extra_3_1_ruser_data -> tg3_1:ruser_data
	wire    [3:0] tg3_1_axi_extra_wuser_strb;                       // tg3_1:wuser_strb -> hbm_0_example_design:axi_extra_3_1_wuser_strb
	wire   [31:0] tg3_1_axi_extra_wuser_data;                       // tg3_1:wuser_data -> hbm_0_example_design:axi_extra_3_1_wuser_data
	wire          hbm_0_example_design_axi_extra_4_0_ruser_err_dbe; // hbm_0_example_design:axi_extra_4_0_ruser_err_dbe -> tg4_0:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_4_0_ruser_data;    // hbm_0_example_design:axi_extra_4_0_ruser_data -> tg4_0:ruser_data
	wire    [3:0] tg4_0_axi_extra_wuser_strb;                       // tg4_0:wuser_strb -> hbm_0_example_design:axi_extra_4_0_wuser_strb
	wire   [31:0] tg4_0_axi_extra_wuser_data;                       // tg4_0:wuser_data -> hbm_0_example_design:axi_extra_4_0_wuser_data
	wire          hbm_0_example_design_axi_extra_4_1_ruser_err_dbe; // hbm_0_example_design:axi_extra_4_1_ruser_err_dbe -> tg4_1:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_4_1_ruser_data;    // hbm_0_example_design:axi_extra_4_1_ruser_data -> tg4_1:ruser_data
	wire    [3:0] tg4_1_axi_extra_wuser_strb;                       // tg4_1:wuser_strb -> hbm_0_example_design:axi_extra_4_1_wuser_strb
	wire   [31:0] tg4_1_axi_extra_wuser_data;                       // tg4_1:wuser_data -> hbm_0_example_design:axi_extra_4_1_wuser_data
	wire          hbm_0_example_design_axi_extra_5_0_ruser_err_dbe; // hbm_0_example_design:axi_extra_5_0_ruser_err_dbe -> tg5_0:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_5_0_ruser_data;    // hbm_0_example_design:axi_extra_5_0_ruser_data -> tg5_0:ruser_data
	wire    [3:0] tg5_0_axi_extra_wuser_strb;                       // tg5_0:wuser_strb -> hbm_0_example_design:axi_extra_5_0_wuser_strb
	wire   [31:0] tg5_0_axi_extra_wuser_data;                       // tg5_0:wuser_data -> hbm_0_example_design:axi_extra_5_0_wuser_data
	wire          hbm_0_example_design_axi_extra_5_1_ruser_err_dbe; // hbm_0_example_design:axi_extra_5_1_ruser_err_dbe -> tg5_1:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_5_1_ruser_data;    // hbm_0_example_design:axi_extra_5_1_ruser_data -> tg5_1:ruser_data
	wire    [3:0] tg5_1_axi_extra_wuser_strb;                       // tg5_1:wuser_strb -> hbm_0_example_design:axi_extra_5_1_wuser_strb
	wire   [31:0] tg5_1_axi_extra_wuser_data;                       // tg5_1:wuser_data -> hbm_0_example_design:axi_extra_5_1_wuser_data
	wire          hbm_0_example_design_axi_extra_6_0_ruser_err_dbe; // hbm_0_example_design:axi_extra_6_0_ruser_err_dbe -> tg6_0:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_6_0_ruser_data;    // hbm_0_example_design:axi_extra_6_0_ruser_data -> tg6_0:ruser_data
	wire    [3:0] tg6_0_axi_extra_wuser_strb;                       // tg6_0:wuser_strb -> hbm_0_example_design:axi_extra_6_0_wuser_strb
	wire   [31:0] tg6_0_axi_extra_wuser_data;                       // tg6_0:wuser_data -> hbm_0_example_design:axi_extra_6_0_wuser_data
	wire          hbm_0_example_design_axi_extra_6_1_ruser_err_dbe; // hbm_0_example_design:axi_extra_6_1_ruser_err_dbe -> tg6_1:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_6_1_ruser_data;    // hbm_0_example_design:axi_extra_6_1_ruser_data -> tg6_1:ruser_data
	wire    [3:0] tg6_1_axi_extra_wuser_strb;                       // tg6_1:wuser_strb -> hbm_0_example_design:axi_extra_6_1_wuser_strb
	wire   [31:0] tg6_1_axi_extra_wuser_data;                       // tg6_1:wuser_data -> hbm_0_example_design:axi_extra_6_1_wuser_data
	wire          hbm_0_example_design_axi_extra_7_0_ruser_err_dbe; // hbm_0_example_design:axi_extra_7_0_ruser_err_dbe -> tg7_0:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_7_0_ruser_data;    // hbm_0_example_design:axi_extra_7_0_ruser_data -> tg7_0:ruser_data
	wire    [3:0] tg7_0_axi_extra_wuser_strb;                       // tg7_0:wuser_strb -> hbm_0_example_design:axi_extra_7_0_wuser_strb
	wire   [31:0] tg7_0_axi_extra_wuser_data;                       // tg7_0:wuser_data -> hbm_0_example_design:axi_extra_7_0_wuser_data
	wire          hbm_0_example_design_axi_extra_7_1_ruser_err_dbe; // hbm_0_example_design:axi_extra_7_1_ruser_err_dbe -> tg7_1:ruser_err_dbe
	wire   [31:0] hbm_0_example_design_axi_extra_7_1_ruser_data;    // hbm_0_example_design:axi_extra_7_1_ruser_data -> tg7_1:ruser_data
	wire    [3:0] tg7_1_axi_extra_wuser_strb;                       // tg7_1:wuser_strb -> hbm_0_example_design:axi_extra_7_1_wuser_strb
	wire   [31:0] tg7_1_axi_extra_wuser_data;                       // tg7_1:wuser_data -> hbm_0_example_design:axi_extra_7_1_wuser_data
	wire          core_clk_iopll_locked_export;                     // core_clk_iopll:locked -> hbm_0_example_design:ext_core_clk_locked
	wire          reset_release_ip_ninit_done_ninit_done;           // reset_release_ip:ninit_done -> ninit_done_splitter:sig_input
	wire          ninit_done_splitter_sig_output_if_0_ninit_done;   // ninit_done_splitter:sig_output_0 -> tg0_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_1_ninit_done;   // ninit_done_splitter:sig_output_1 -> tg0_1:ninit_done
	wire          ninit_done_splitter_sig_output_if_10_ninit_done;  // ninit_done_splitter:sig_output_10 -> tg5_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_11_ninit_done;  // ninit_done_splitter:sig_output_11 -> tg5_1:ninit_done
	wire          ninit_done_splitter_sig_output_if_12_ninit_done;  // ninit_done_splitter:sig_output_12 -> tg6_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_13_ninit_done;  // ninit_done_splitter:sig_output_13 -> tg6_1:ninit_done
	wire          ninit_done_splitter_sig_output_if_14_ninit_done;  // ninit_done_splitter:sig_output_14 -> tg7_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_15_ninit_done;  // ninit_done_splitter:sig_output_15 -> tg7_1:ninit_done
	wire          ninit_done_splitter_sig_output_if_2_ninit_done;   // ninit_done_splitter:sig_output_2 -> tg1_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_3_ninit_done;   // ninit_done_splitter:sig_output_3 -> tg1_1:ninit_done
	wire          ninit_done_splitter_sig_output_if_4_ninit_done;   // ninit_done_splitter:sig_output_4 -> tg2_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_5_ninit_done;   // ninit_done_splitter:sig_output_5 -> tg2_1:ninit_done
	wire          ninit_done_splitter_sig_output_if_6_ninit_done;   // ninit_done_splitter:sig_output_6 -> tg3_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_7_ninit_done;   // ninit_done_splitter:sig_output_7 -> tg3_1:ninit_done
	wire          ninit_done_splitter_sig_output_if_8_ninit_done;   // ninit_done_splitter:sig_output_8 -> tg4_0:ninit_done
	wire          ninit_done_splitter_sig_output_if_9_ninit_done;   // ninit_done_splitter:sig_output_9 -> tg4_1:ninit_done
	wire          hbm_0_example_design_wmcrst_n_0_reset;            // hbm_0_example_design:wmcrst_n_0 -> [tg0_0:wmcrst_n_in, tg0_1:wmcrst_n_in, tg1_0:wmcrst_n_in, tg1_1:wmcrst_n_in]
	wire          hbm_0_example_design_wmcrst_n_2_reset;            // hbm_0_example_design:wmcrst_n_2 -> [tg2_0:wmcrst_n_in, tg2_1:wmcrst_n_in, tg3_0:wmcrst_n_in, tg3_1:wmcrst_n_in]
	wire          hbm_0_example_design_wmcrst_n_4_reset;            // hbm_0_example_design:wmcrst_n_4 -> [tg4_0:wmcrst_n_in, tg4_1:wmcrst_n_in, tg5_0:wmcrst_n_in, tg5_1:wmcrst_n_in]
	wire          hbm_0_example_design_wmcrst_n_6_reset;            // hbm_0_example_design:wmcrst_n_6 -> [tg6_0:wmcrst_n_in, tg6_1:wmcrst_n_in, tg7_0:wmcrst_n_in, tg7_1:wmcrst_n_in]

  //-- axi slave signals {{{
  wire [13:0] s0_awaddr;
  wire [2:0] s0_awprot;
  wire s0_awvalid;
  wire s0_awready;

  wire [31:0] s0_wdata;
  wire [3:0] s0_wstrb;
  wire s0_wvalid;
  wire s0_wready;

  wire [1:0] s0_bresp;
  wire s0_bvalid;
  wire s0_bready;

  wire [13:0] s0_araddr;
  wire [2:0] s0_arprot;
  wire s0_arvalid;
  wire s0_arready;

  wire [31:0] s0_rdata;
  wire [1:0] s0_rresp;
  wire s0_rvalid;
  wire s0_rready;
  //-- axi master wires {{{
  //-- interface 0 {{{
  //-- ar channel
  wire [31:0] m0_araddr;
  wire [7:0] m0_arlen;
  wire [2:0] m0_arsize;
  wire [1:0] m0_arburst;
  wire m0_arvalid;
  wire m0_arready;
  wire [6:0] m0_arid;
  //-- r channel
  wire [1023:0] m0_rdata;
  wire [1:0] m0_rresp;
  wire m0_rlast;
  wire m0_rvalid;
  wire m0_rready;
  wire [6:0] m0_rid;
  //-- aw channel
  wire [31:0] m0_awaddr ;
  wire m0_awvalid;
  wire m0_awready;
  wire [7:0] m0_awlen;
  wire [2:0] m0_awsize;
  wire [1:0] m0_awburst;
  wire [6:0] m0_awid;
  //-- w channel
  wire [1023:0] m0_wdata;
  wire [127:0] m0_wstrb;
  wire m0_wlast;
  wire m0_wvalid;
  wire m0_wready;
  //-- b channel
  wire m0_bvalid;
  wire m0_bready;
  wire [6:0] m0_bid;
  //--}}}
  //-- interface 1 {{{
  //-- ar channel
  wire [31:0] m1_araddr;
  wire [7:0] m1_arlen;
  wire [2:0] m1_arsize;
  wire [1:0] m1_arburst;
  wire m1_arvalid;
  wire m1_arready;
  wire [6:0] m1_arid;
  //-- r channel
  wire [1023:0] m1_rdata;
  wire [1:0] m1_rresp;
  wire m1_rlast;
  wire m1_rvalid;
  wire m1_rready;
  wire [6:0] m1_rid;
  //-- aw channel
  wire [31:0] m1_awaddr;
  wire m1_awvalid;
  wire m1_awready;
  wire [7:0] m1_awlen;
  wire [2:0] m1_awsize;
  wire [1:0] m1_awburst;
  wire [6:0] m1_awid;
  //-- w channel
  wire [1023:0] m1_wdata;
  wire [127:0] m1_wstrb;
  wire m1_wlast;
  wire m1_wvalid;
  wire m1_wready;
  //-- b channel
  wire m1_bvalid;
  wire m1_bready;
  wire [6:0] m1_bid;
  //--}}}
  //-- interface 2 {{{
  //-- ar channel
  wire [31:0] m2_araddr;
  wire [7:0] m2_arlen;
  wire [2:0] m2_arsize;
  wire [1:0] m2_arburst;
  wire m2_arvalid;
  wire m2_arready;
  wire [6:0] m2_arid;
  //-- r channel
  wire [1023:0] m2_rdata;
  wire [1:0] m2_rresp;
  wire m2_rlast;
  wire m2_rvalid;
  wire m2_rready;
  wire [6:0] m2_rid;
  //-- aw channel
  wire [31:0] m2_awaddr;
  wire m2_awvalid;
  wire m2_awready;
  wire [7:0] m2_awlen;
  wire [2:0] m2_awsize;
  wire [1:0] m2_awburst;
  wire [6:0] m2_awid;
  //-- w channel
  wire [1023:0] m2_wdata;
  wire [127:0] m2_wstrb;
  wire m2_wlast;
  wire m2_wvalid;
  wire m2_wready;
  //-- b channel
  wire m2_bvalid;
  wire m2_bready;
  wire [6:0] m2_bid;
  //--}}}
  //-- interface 3 {{{
  //-- ar channel
  wire [31:0] m3_araddr;
  wire [7:0] m3_arlen;
  wire [2:0] m3_arsize;
  wire [1:0] m3_arburst;
  wire m3_arvalid;
  wire m3_arready;
  wire [6:0] m3_arid;
  //-- r channel
  wire [1023:0] m3_rdata;
  wire [1:0] m3_rresp;
  wire m3_rlast;
  wire m3_rvalid;
  wire m3_rready;
  wire [6:0] m3_rid;
  //-- aw channel
  wire [31:0] m3_awaddr;
  wire m3_awvalid;
  wire m3_awready;
  wire [7:0] m3_awlen;
  wire [2:0] m3_awsize;
  wire [1:0] m3_awburst;
  wire [6:0] m3_awid;
  //-- w channel
  wire [1023:0] m3_wdata;
  wire [127:0] m3_wstrb;
  wire m3_wlast;
  wire m3_wvalid;
  wire m3_wready;
  //-- b channel
  wire m3_bvalid;
  wire m3_bready;
  wire [6:0] m3_bid;

	ed_synth_core_clk_iopll core_clk_iopll (
		.rst      (core_clk_iopll_reset_reset),   //   input,  width = 1,   reset.reset
		.refclk   (core_clk_iopll_ref_clk_clk),   //   input,  width = 1,  refclk.clk
		.locked   (core_clk_iopll_locked_export), //  output,  width = 1,  locked.export
		.outclk_0 (core_clk_iopll_outclk0_clk)    //  output,  width = 1, outclk0.clk
	);

	ed_synth_hbm_0_example_design hbm_0_example_design (
		.pll_ref_clk                 (hbm_0_example_design_pll_ref_clk_clk),             //   input,    width = 1,         pll_ref_clk.clk
		.ext_core_clk                (core_clk_iopll_outclk0_clk),                       //   input,    width = 1,        ext_core_clk.clk
		.ext_core_clk_locked         (core_clk_iopll_locked_export),                     //   input,    width = 1, ext_core_clk_locked.export
		.wmcrst_n_in                 (hbm_0_example_design_wmcrst_n_in_reset_n),         //   input,    width = 1,         wmcrst_n_in.reset_n
		.hbm_only_reset_in           (hbm_only_reset_in_reset),                          //   input,    width = 1,   hbm_only_reset_in.reset
		.local_cal_success           (),                                                 //  output,    width = 1,              status.local_cal_success
		.local_cal_fail              (),                                                 //  output,    width = 1,                    .local_cal_fail
		.cal_lat                     (),                                                 //  output,    width = 3,             cal_lat.cal_lat
		.ck_t_0                      (),                                                 //  output,    width = 1,               mem_0.ck_t
		.ck_c_0                      (),                                                 //  output,    width = 1,                    .ck_c
		.cke_0                       (),                                                 //  output,    width = 1,                    .cke
		.c_0                         (),                                                 //  output,    width = 8,                    .c
		.r_0                         (),                                                 //  output,    width = 6,                    .r
		.dq_0                        (),                                                 //   inout,  width = 128,                    .dq
		.dm_0                        (),                                                 //   inout,   width = 16,                    .dm
		.dbi_0                       (),                                                 //   inout,   width = 16,                    .dbi
		.par_0                       (),                                                 //   inout,    width = 4,                    .par
		.derr_0                      (),                                                 //   inout,    width = 4,                    .derr
		.rdqs_t_0                    (),                                                 //   input,    width = 4,                    .rdqs_t
		.rdqs_c_0                    (),                                                 //   input,    width = 4,                    .rdqs_c
		.wdqs_t_0                    (),                                                 //  output,    width = 4,                    .wdqs_t
		.wdqs_c_0                    (),                                                 //  output,    width = 4,                    .wdqs_c
		.rd_0                        (),                                                 //   inout,    width = 8,                    .rd
		.rr_0                        (),                                                 //  output,    width = 1,                    .rr
		.rc_0                        (),                                                 //  output,    width = 1,                    .rc
		.aerr_0                      (),                                                 //   input,    width = 1,                    .aerr
		.ck_t_1                      (),                                                 //  output,    width = 1,               mem_1.ck_t
		.ck_c_1                      (),                                                 //  output,    width = 1,                    .ck_c
		.cke_1                       (),                                                 //  output,    width = 1,                    .cke
		.c_1                         (),                                                 //  output,    width = 8,                    .c
		.r_1                         (),                                                 //  output,    width = 6,                    .r
		.dq_1                        (),                                                 //   inout,  width = 128,                    .dq
		.dm_1                        (),                                                 //   inout,   width = 16,                    .dm
		.dbi_1                       (),                                                 //   inout,   width = 16,                    .dbi
		.par_1                       (),                                                 //   inout,    width = 4,                    .par
		.derr_1                      (),                                                 //   inout,    width = 4,                    .derr
		.rdqs_t_1                    (),                                                 //   input,    width = 4,                    .rdqs_t
		.rdqs_c_1                    (),                                                 //   input,    width = 4,                    .rdqs_c
		.wdqs_t_1                    (),                                                 //  output,    width = 4,                    .wdqs_t
		.wdqs_c_1                    (),                                                 //  output,    width = 4,                    .wdqs_c
		.rd_1                        (),                                                 //   inout,    width = 8,                    .rd
		.rr_1                        (),                                                 //  output,    width = 1,                    .rr
		.rc_1                        (),                                                 //  output,    width = 1,                    .rc
		.aerr_1                      (),                                                 //   input,    width = 1,                    .aerr
		.ck_t_2                      (),                                                 //  output,    width = 1,               mem_2.ck_t
		.ck_c_2                      (),                                                 //  output,    width = 1,                    .ck_c
		.cke_2                       (),                                                 //  output,    width = 1,                    .cke
		.c_2                         (),                                                 //  output,    width = 8,                    .c
		.r_2                         (),                                                 //  output,    width = 6,                    .r
		.dq_2                        (),                                                 //   inout,  width = 128,                    .dq
		.dm_2                        (),                                                 //   inout,   width = 16,                    .dm
		.dbi_2                       (),                                                 //   inout,   width = 16,                    .dbi
		.par_2                       (),                                                 //   inout,    width = 4,                    .par
		.derr_2                      (),                                                 //   inout,    width = 4,                    .derr
		.rdqs_t_2                    (),                                                 //   input,    width = 4,                    .rdqs_t
		.rdqs_c_2                    (),                                                 //   input,    width = 4,                    .rdqs_c
		.wdqs_t_2                    (),                                                 //  output,    width = 4,                    .wdqs_t
		.wdqs_c_2                    (),                                                 //  output,    width = 4,                    .wdqs_c
		.rd_2                        (),                                                 //   inout,    width = 8,                    .rd
		.rr_2                        (),                                                 //  output,    width = 1,                    .rr
		.rc_2                        (),                                                 //  output,    width = 1,                    .rc
		.aerr_2                      (),                                                 //   input,    width = 1,                    .aerr
		.ck_t_3                      (),                                                 //  output,    width = 1,               mem_3.ck_t
		.ck_c_3                      (),                                                 //  output,    width = 1,                    .ck_c
		.cke_3                       (),                                                 //  output,    width = 1,                    .cke
		.c_3                         (),                                                 //  output,    width = 8,                    .c
		.r_3                         (),                                                 //  output,    width = 6,                    .r
		.dq_3                        (),                                                 //   inout,  width = 128,                    .dq
		.dm_3                        (),                                                 //   inout,   width = 16,                    .dm
		.dbi_3                       (),                                                 //   inout,   width = 16,                    .dbi
		.par_3                       (),                                                 //   inout,    width = 4,                    .par
		.derr_3                      (),                                                 //   inout,    width = 4,                    .derr
		.rdqs_t_3                    (),                                                 //   input,    width = 4,                    .rdqs_t
		.rdqs_c_3                    (),                                                 //   input,    width = 4,                    .rdqs_c
		.wdqs_t_3                    (),                                                 //  output,    width = 4,                    .wdqs_t
		.wdqs_c_3                    (),                                                 //  output,    width = 4,                    .wdqs_c
		.rd_3                        (),                                                 //   inout,    width = 8,                    .rd
		.rr_3                        (),                                                 //  output,    width = 1,                    .rr
		.rc_3                        (),                                                 //  output,    width = 1,                    .rc
		.aerr_3                      (),                                                 //   input,    width = 1,                    .aerr
		.ck_t_4                      (),                                                 //  output,    width = 1,               mem_4.ck_t
		.ck_c_4                      (),                                                 //  output,    width = 1,                    .ck_c
		.cke_4                       (),                                                 //  output,    width = 1,                    .cke
		.c_4                         (),                                                 //  output,    width = 8,                    .c
		.r_4                         (),                                                 //  output,    width = 6,                    .r
		.dq_4                        (),                                                 //   inout,  width = 128,                    .dq
		.dm_4                        (),                                                 //   inout,   width = 16,                    .dm
		.dbi_4                       (),                                                 //   inout,   width = 16,                    .dbi
		.par_4                       (),                                                 //   inout,    width = 4,                    .par
		.derr_4                      (),                                                 //   inout,    width = 4,                    .derr
		.rdqs_t_4                    (),                                                 //   input,    width = 4,                    .rdqs_t
		.rdqs_c_4                    (),                                                 //   input,    width = 4,                    .rdqs_c
		.wdqs_t_4                    (),                                                 //  output,    width = 4,                    .wdqs_t
		.wdqs_c_4                    (),                                                 //  output,    width = 4,                    .wdqs_c
		.rd_4                        (),                                                 //   inout,    width = 8,                    .rd
		.rr_4                        (),                                                 //  output,    width = 1,                    .rr
		.rc_4                        (),                                                 //  output,    width = 1,                    .rc
		.aerr_4                      (),                                                 //   input,    width = 1,                    .aerr
		.ck_t_5                      (),                                                 //  output,    width = 1,               mem_5.ck_t
		.ck_c_5                      (),                                                 //  output,    width = 1,                    .ck_c
		.cke_5                       (),                                                 //  output,    width = 1,                    .cke
		.c_5                         (),                                                 //  output,    width = 8,                    .c
		.r_5                         (),                                                 //  output,    width = 6,                    .r
		.dq_5                        (),                                                 //   inout,  width = 128,                    .dq
		.dm_5                        (),                                                 //   inout,   width = 16,                    .dm
		.dbi_5                       (),                                                 //   inout,   width = 16,                    .dbi
		.par_5                       (),                                                 //   inout,    width = 4,                    .par
		.derr_5                      (),                                                 //   inout,    width = 4,                    .derr
		.rdqs_t_5                    (),                                                 //   input,    width = 4,                    .rdqs_t
		.rdqs_c_5                    (),                                                 //   input,    width = 4,                    .rdqs_c
		.wdqs_t_5                    (),                                                 //  output,    width = 4,                    .wdqs_t
		.wdqs_c_5                    (),                                                 //  output,    width = 4,                    .wdqs_c
		.rd_5                        (),                                                 //   inout,    width = 8,                    .rd
		.rr_5                        (),                                                 //  output,    width = 1,                    .rr
		.rc_5                        (),                                                 //  output,    width = 1,                    .rc
		.aerr_5                      (),                                                 //   input,    width = 1,                    .aerr
		.ck_t_6                      (),                                                 //  output,    width = 1,               mem_6.ck_t
		.ck_c_6                      (),                                                 //  output,    width = 1,                    .ck_c
		.cke_6                       (),                                                 //  output,    width = 1,                    .cke
		.c_6                         (),                                                 //  output,    width = 8,                    .c
		.r_6                         (),                                                 //  output,    width = 6,                    .r
		.dq_6                        (),                                                 //   inout,  width = 128,                    .dq
		.dm_6                        (),                                                 //   inout,   width = 16,                    .dm
		.dbi_6                       (),                                                 //   inout,   width = 16,                    .dbi
		.par_6                       (),                                                 //   inout,    width = 4,                    .par
		.derr_6                      (),                                                 //   inout,    width = 4,                    .derr
		.rdqs_t_6                    (),                                                 //   input,    width = 4,                    .rdqs_t
		.rdqs_c_6                    (),                                                 //   input,    width = 4,                    .rdqs_c
		.wdqs_t_6                    (),                                                 //  output,    width = 4,                    .wdqs_t
		.wdqs_c_6                    (),                                                 //  output,    width = 4,                    .wdqs_c
		.rd_6                        (),                                                 //   inout,    width = 8,                    .rd
		.rr_6                        (),                                                 //  output,    width = 1,                    .rr
		.rc_6                        (),                                                 //  output,    width = 1,                    .rc
		.aerr_6                      (),                                                 //   input,    width = 1,                    .aerr
		.ck_t_7                      (),                                                 //  output,    width = 1,               mem_7.ck_t
		.ck_c_7                      (),                                                 //  output,    width = 1,                    .ck_c
		.cke_7                       (),                                                 //  output,    width = 1,                    .cke
		.c_7                         (),                                                 //  output,    width = 8,                    .c
		.r_7                         (),                                                 //  output,    width = 6,                    .r
		.dq_7                        (),                                                 //   inout,  width = 128,                    .dq
		.dm_7                        (),                                                 //   inout,   width = 16,                    .dm
		.dbi_7                       (),                                                 //   inout,   width = 16,                    .dbi
		.par_7                       (),                                                 //   inout,    width = 4,                    .par
		.derr_7                      (),                                                 //   inout,    width = 4,                    .derr
		.rdqs_t_7                    (),                                                 //   input,    width = 4,                    .rdqs_t
		.rdqs_c_7                    (),                                                 //   input,    width = 4,                    .rdqs_c
		.wdqs_t_7                    (),                                                 //  output,    width = 4,                    .wdqs_t
		.wdqs_c_7                    (),                                                 //  output,    width = 4,                    .wdqs_c
		.rd_7                        (),                                                 //   inout,    width = 8,                    .rd
		.rr_7                        (),                                                 //  output,    width = 1,                    .rr
		.rc_7                        (),                                                 //  output,    width = 1,                    .rc
		.aerr_7                      (),                                                 //   input,    width = 1,                    .aerr
		.cattrip                     (m2u_bridge_cattrip),                               //   input,    width = 1,          m2u_bridge.cattrip
		.temp                        (m2u_bridge_temp),                                  //   input,    width = 3,                    .temp
		.wso                         (m2u_bridge_wso),                                   //   input,    width = 8,                    .wso
		.reset_n                     (m2u_bridge_reset_n),                               //  output,    width = 1,                    .reset_n
		.wrst_n                      (m2u_bridge_wrst_n),                                //  output,    width = 1,                    .wrst_n
		.wrck                        (m2u_bridge_wrck),                                  //  output,    width = 1,                    .wrck
		.shiftwr                     (m2u_bridge_shiftwr),                               //  output,    width = 1,                    .shiftwr
		.capturewr                   (m2u_bridge_capturewr),                             //  output,    width = 1,                    .capturewr
		.updatewr                    (m2u_bridge_updatewr),                              //  output,    width = 1,                    .updatewr
		.selectwir                   (m2u_bridge_selectwir),                             //  output,    width = 1,                    .selectwir
		.wsi                         (m2u_bridge_wsi),                                   //  output,    width = 1,                    .wsi
		.phy_clk_0_clk               (),                                                 //  output,    width = 1,           phy_clk_0.clk
		.axi_extra_0_0_ruser_err_dbe (hbm_0_example_design_axi_extra_0_0_ruser_err_dbe), //  output,    width = 1,       axi_extra_0_0.ruser_err_dbe
		.axi_extra_0_0_ruser_data    (hbm_0_example_design_axi_extra_0_0_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_0_0_wuser_data    (tg0_0_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_0_0_wuser_strb    (tg0_0_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_0_1_ruser_err_dbe (hbm_0_example_design_axi_extra_0_1_ruser_err_dbe), //  output,    width = 1,       axi_extra_0_1.ruser_err_dbe
		.axi_extra_0_1_ruser_data    (hbm_0_example_design_axi_extra_0_1_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_0_1_wuser_data    (tg0_1_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_0_1_wuser_strb    (tg0_1_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_1_0_ruser_err_dbe (hbm_0_example_design_axi_extra_1_0_ruser_err_dbe), //  output,    width = 1,       axi_extra_1_0.ruser_err_dbe
		.axi_extra_1_0_ruser_data    (hbm_0_example_design_axi_extra_1_0_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_1_0_wuser_data    (tg1_0_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_1_0_wuser_strb    (tg1_0_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_1_1_ruser_err_dbe (hbm_0_example_design_axi_extra_1_1_ruser_err_dbe), //  output,    width = 1,       axi_extra_1_1.ruser_err_dbe
		.axi_extra_1_1_ruser_data    (hbm_0_example_design_axi_extra_1_1_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_1_1_wuser_data    (tg1_1_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_1_1_wuser_strb    (tg1_1_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.apb_0_ur_paddr              (tg0_0_apb_ur_paddr),                               //   input,   width = 16,               apb_0.ur_paddr
		.apb_0_ur_psel               (tg0_0_apb_ur_psel),                                //   input,    width = 1,                    .ur_psel
		.apb_0_ur_penable            (tg0_0_apb_ur_penable),                             //   input,    width = 1,                    .ur_penable
		.apb_0_ur_pwrite             (tg0_0_apb_ur_pwrite),                              //   input,    width = 1,                    .ur_pwrite
		.apb_0_ur_pwdata             (tg0_0_apb_ur_pwdata),                              //   input,   width = 16,                    .ur_pwdata
		.apb_0_ur_pstrb              (tg0_0_apb_ur_pstrb),                               //   input,    width = 2,                    .ur_pstrb
		.apb_0_ur_prready            (hbm_0_example_design_apb_0_ur_prready),            //  output,    width = 1,                    .ur_prready
		.apb_0_ur_prdata             (hbm_0_example_design_apb_0_ur_prdata),             //  output,   width = 16,                    .ur_prdata
		.apb_1_ur_paddr              (tg1_0_apb_ur_paddr),                               //   input,   width = 16,               apb_1.ur_paddr
		.apb_1_ur_psel               (tg1_0_apb_ur_psel),                                //   input,    width = 1,                    .ur_psel
		.apb_1_ur_penable            (tg1_0_apb_ur_penable),                             //   input,    width = 1,                    .ur_penable
		.apb_1_ur_pwrite             (tg1_0_apb_ur_pwrite),                              //   input,    width = 1,                    .ur_pwrite
		.apb_1_ur_pwdata             (tg1_0_apb_ur_pwdata),                              //   input,   width = 16,                    .ur_pwdata
		.apb_1_ur_pstrb              (tg1_0_apb_ur_pstrb),                               //   input,    width = 2,                    .ur_pstrb
		.apb_1_ur_prready            (hbm_0_example_design_apb_1_ur_prready),            //  output,    width = 1,                    .ur_prready
		.apb_1_ur_prdata             (hbm_0_example_design_apb_1_ur_prdata),             //  output,   width = 16,                    .ur_prdata
		.axi_0_0_awid                (tg0_0_axi_awid),                                   //   input,    width = 7,             axi_0_0.awid
		.axi_0_0_awaddr              (tg0_0_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_0_0_awlen               (tg0_0_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_0_0_awsize              (tg0_0_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_0_0_awburst             (tg0_0_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_0_0_awprot              (tg0_0_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_0_0_awqos               (tg0_0_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_0_0_awuser              (tg0_0_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_0_0_awvalid             (tg0_0_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_0_0_awready             (tg0_0_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_0_0_wdata               (tg0_0_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_0_0_wstrb               (tg0_0_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_0_0_wlast               (tg0_0_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_0_0_wvalid              (tg0_0_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_0_0_wready              (tg0_0_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_0_0_bid                 (tg0_0_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_0_0_bresp               (tg0_0_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_0_0_bvalid              (tg0_0_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_0_0_bready              (tg0_0_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_0_0_arid                (tg0_0_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_0_0_araddr              (tg0_0_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_0_0_arlen               (tg0_0_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_0_0_arsize              (tg0_0_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_0_0_arburst             (tg0_0_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_0_0_arprot              (tg0_0_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_0_0_arqos               (tg0_0_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_0_0_aruser              (tg0_0_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_0_0_arvalid             (tg0_0_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_0_0_arready             (tg0_0_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_0_0_rid                 (tg0_0_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_0_0_rdata               (tg0_0_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_0_0_rresp               (tg0_0_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_0_0_rlast               (tg0_0_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_0_0_rvalid              (tg0_0_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_0_0_rready              (tg0_0_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_0_1_awid                (tg0_1_axi_awid),                                   //   input,    width = 7,             axi_0_1.awid
		.axi_0_1_awaddr              (tg0_1_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_0_1_awlen               (tg0_1_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_0_1_awsize              (tg0_1_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_0_1_awburst             (tg0_1_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_0_1_awprot              (tg0_1_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_0_1_awqos               (tg0_1_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_0_1_awuser              (tg0_1_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_0_1_awvalid             (tg0_1_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_0_1_awready             (tg0_1_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_0_1_wdata               (tg0_1_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_0_1_wstrb               (tg0_1_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_0_1_wlast               (tg0_1_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_0_1_wvalid              (tg0_1_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_0_1_wready              (tg0_1_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_0_1_bid                 (tg0_1_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_0_1_bresp               (tg0_1_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_0_1_bvalid              (tg0_1_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_0_1_bready              (tg0_1_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_0_1_arid                (tg0_1_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_0_1_araddr              (tg0_1_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_0_1_arlen               (tg0_1_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_0_1_arsize              (tg0_1_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_0_1_arburst             (tg0_1_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_0_1_arprot              (tg0_1_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_0_1_arqos               (tg0_1_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_0_1_aruser              (tg0_1_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_0_1_arvalid             (tg0_1_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_0_1_arready             (tg0_1_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_0_1_rid                 (tg0_1_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_0_1_rdata               (tg0_1_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_0_1_rresp               (tg0_1_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_0_1_rlast               (tg0_1_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_0_1_rvalid              (tg0_1_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_0_1_rready              (tg0_1_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_1_0_awid                (tg1_0_axi_awid),                                   //   input,    width = 7,             axi_1_0.awid
		.axi_1_0_awaddr              (tg1_0_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_1_0_awlen               (tg1_0_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_1_0_awsize              (tg1_0_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_1_0_awburst             (tg1_0_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_1_0_awprot              (tg1_0_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_1_0_awqos               (tg1_0_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_1_0_awuser              (tg1_0_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_1_0_awvalid             (tg1_0_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_1_0_awready             (tg1_0_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_1_0_wdata               (tg1_0_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_1_0_wstrb               (tg1_0_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_1_0_wlast               (tg1_0_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_1_0_wvalid              (tg1_0_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_1_0_wready              (tg1_0_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_1_0_bid                 (tg1_0_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_1_0_bresp               (tg1_0_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_1_0_bvalid              (tg1_0_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_1_0_bready              (tg1_0_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_1_0_arid                (tg1_0_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_1_0_araddr              (tg1_0_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_1_0_arlen               (tg1_0_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_1_0_arsize              (tg1_0_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_1_0_arburst             (tg1_0_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_1_0_arprot              (tg1_0_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_1_0_arqos               (tg1_0_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_1_0_aruser              (tg1_0_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_1_0_arvalid             (tg1_0_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_1_0_arready             (tg1_0_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_1_0_rid                 (tg1_0_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_1_0_rdata               (tg1_0_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_1_0_rresp               (tg1_0_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_1_0_rlast               (tg1_0_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_1_0_rvalid              (tg1_0_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_1_0_rready              (tg1_0_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_1_1_awid                (tg1_1_axi_awid),                                   //   input,    width = 7,             axi_1_1.awid
		.axi_1_1_awaddr              (tg1_1_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_1_1_awlen               (tg1_1_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_1_1_awsize              (tg1_1_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_1_1_awburst             (tg1_1_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_1_1_awprot              (tg1_1_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_1_1_awqos               (tg1_1_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_1_1_awuser              (tg1_1_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_1_1_awvalid             (tg1_1_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_1_1_awready             (tg1_1_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_1_1_wdata               (tg1_1_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_1_1_wstrb               (tg1_1_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_1_1_wlast               (tg1_1_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_1_1_wvalid              (tg1_1_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_1_1_wready              (tg1_1_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_1_1_bid                 (tg1_1_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_1_1_bresp               (tg1_1_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_1_1_bvalid              (tg1_1_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_1_1_bready              (tg1_1_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_1_1_arid                (tg1_1_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_1_1_araddr              (tg1_1_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_1_1_arlen               (tg1_1_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_1_1_arsize              (tg1_1_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_1_1_arburst             (tg1_1_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_1_1_arprot              (tg1_1_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_1_1_arqos               (tg1_1_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_1_1_aruser              (tg1_1_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_1_1_arvalid             (tg1_1_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_1_1_arready             (tg1_1_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_1_1_rid                 (tg1_1_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_1_1_rdata               (tg1_1_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_1_1_rresp               (tg1_1_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_1_1_rlast               (tg1_1_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_1_1_rvalid              (tg1_1_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_1_1_rready              (tg1_1_axi_rready),                                 //   input,    width = 1,                    .rready
		.wmc_clk_0                   (hbm_0_example_design_wmc_clk_0_clk),               //  output,    width = 1,           wmc_clk_0.clk
		.wmcrst_n_0                  (hbm_0_example_design_wmcrst_n_0_reset),            //  output,    width = 1,          wmcrst_n_0.reset_n
		.phy_clk_2_clk               (),                                                 //  output,    width = 1,           phy_clk_2.clk
		.axi_extra_2_0_ruser_err_dbe (hbm_0_example_design_axi_extra_2_0_ruser_err_dbe), //  output,    width = 1,       axi_extra_2_0.ruser_err_dbe
		.axi_extra_2_0_ruser_data    (hbm_0_example_design_axi_extra_2_0_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_2_0_wuser_data    (tg2_0_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_2_0_wuser_strb    (tg2_0_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_2_1_ruser_err_dbe (hbm_0_example_design_axi_extra_2_1_ruser_err_dbe), //  output,    width = 1,       axi_extra_2_1.ruser_err_dbe
		.axi_extra_2_1_ruser_data    (hbm_0_example_design_axi_extra_2_1_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_2_1_wuser_data    (tg2_1_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_2_1_wuser_strb    (tg2_1_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_3_0_ruser_err_dbe (hbm_0_example_design_axi_extra_3_0_ruser_err_dbe), //  output,    width = 1,       axi_extra_3_0.ruser_err_dbe
		.axi_extra_3_0_ruser_data    (hbm_0_example_design_axi_extra_3_0_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_3_0_wuser_data    (tg3_0_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_3_0_wuser_strb    (tg3_0_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_3_1_ruser_err_dbe (hbm_0_example_design_axi_extra_3_1_ruser_err_dbe), //  output,    width = 1,       axi_extra_3_1.ruser_err_dbe
		.axi_extra_3_1_ruser_data    (hbm_0_example_design_axi_extra_3_1_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_3_1_wuser_data    (tg3_1_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_3_1_wuser_strb    (tg3_1_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.apb_2_ur_paddr              (tg2_0_apb_ur_paddr),                               //   input,   width = 16,               apb_2.ur_paddr
		.apb_2_ur_psel               (tg2_0_apb_ur_psel),                                //   input,    width = 1,                    .ur_psel
		.apb_2_ur_penable            (tg2_0_apb_ur_penable),                             //   input,    width = 1,                    .ur_penable
		.apb_2_ur_pwrite             (tg2_0_apb_ur_pwrite),                              //   input,    width = 1,                    .ur_pwrite
		.apb_2_ur_pwdata             (tg2_0_apb_ur_pwdata),                              //   input,   width = 16,                    .ur_pwdata
		.apb_2_ur_pstrb              (tg2_0_apb_ur_pstrb),                               //   input,    width = 2,                    .ur_pstrb
		.apb_2_ur_prready            (hbm_0_example_design_apb_2_ur_prready),            //  output,    width = 1,                    .ur_prready
		.apb_2_ur_prdata             (hbm_0_example_design_apb_2_ur_prdata),             //  output,   width = 16,                    .ur_prdata
		.apb_3_ur_paddr              (tg3_0_apb_ur_paddr),                               //   input,   width = 16,               apb_3.ur_paddr
		.apb_3_ur_psel               (tg3_0_apb_ur_psel),                                //   input,    width = 1,                    .ur_psel
		.apb_3_ur_penable            (tg3_0_apb_ur_penable),                             //   input,    width = 1,                    .ur_penable
		.apb_3_ur_pwrite             (tg3_0_apb_ur_pwrite),                              //   input,    width = 1,                    .ur_pwrite
		.apb_3_ur_pwdata             (tg3_0_apb_ur_pwdata),                              //   input,   width = 16,                    .ur_pwdata
		.apb_3_ur_pstrb              (tg3_0_apb_ur_pstrb),                               //   input,    width = 2,                    .ur_pstrb
		.apb_3_ur_prready            (hbm_0_example_design_apb_3_ur_prready),            //  output,    width = 1,                    .ur_prready
		.apb_3_ur_prdata             (hbm_0_example_design_apb_3_ur_prdata),             //  output,   width = 16,                    .ur_prdata
		.axi_2_0_awid                (tg2_0_axi_awid),                                   //   input,    width = 7,             axi_2_0.awid
		.axi_2_0_awaddr              (tg2_0_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_2_0_awlen               (tg2_0_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_2_0_awsize              (tg2_0_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_2_0_awburst             (tg2_0_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_2_0_awprot              (tg2_0_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_2_0_awqos               (tg2_0_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_2_0_awuser              (tg2_0_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_2_0_awvalid             (tg2_0_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_2_0_awready             (tg2_0_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_2_0_wdata               (tg2_0_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_2_0_wstrb               (tg2_0_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_2_0_wlast               (tg2_0_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_2_0_wvalid              (tg2_0_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_2_0_wready              (tg2_0_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_2_0_bid                 (tg2_0_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_2_0_bresp               (tg2_0_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_2_0_bvalid              (tg2_0_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_2_0_bready              (tg2_0_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_2_0_arid                (tg2_0_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_2_0_araddr              (tg2_0_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_2_0_arlen               (tg2_0_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_2_0_arsize              (tg2_0_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_2_0_arburst             (tg2_0_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_2_0_arprot              (tg2_0_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_2_0_arqos               (tg2_0_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_2_0_aruser              (tg2_0_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_2_0_arvalid             (tg2_0_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_2_0_arready             (tg2_0_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_2_0_rid                 (tg2_0_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_2_0_rdata               (tg2_0_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_2_0_rresp               (tg2_0_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_2_0_rlast               (tg2_0_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_2_0_rvalid              (tg2_0_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_2_0_rready              (tg2_0_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_2_1_awid                (tg2_1_axi_awid),                                   //   input,    width = 7,             axi_2_1.awid
		.axi_2_1_awaddr              (tg2_1_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_2_1_awlen               (tg2_1_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_2_1_awsize              (tg2_1_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_2_1_awburst             (tg2_1_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_2_1_awprot              (tg2_1_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_2_1_awqos               (tg2_1_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_2_1_awuser              (tg2_1_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_2_1_awvalid             (tg2_1_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_2_1_awready             (tg2_1_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_2_1_wdata               (tg2_1_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_2_1_wstrb               (tg2_1_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_2_1_wlast               (tg2_1_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_2_1_wvalid              (tg2_1_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_2_1_wready              (tg2_1_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_2_1_bid                 (tg2_1_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_2_1_bresp               (tg2_1_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_2_1_bvalid              (tg2_1_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_2_1_bready              (tg2_1_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_2_1_arid                (tg2_1_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_2_1_araddr              (tg2_1_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_2_1_arlen               (tg2_1_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_2_1_arsize              (tg2_1_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_2_1_arburst             (tg2_1_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_2_1_arprot              (tg2_1_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_2_1_arqos               (tg2_1_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_2_1_aruser              (tg2_1_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_2_1_arvalid             (tg2_1_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_2_1_arready             (tg2_1_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_2_1_rid                 (tg2_1_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_2_1_rdata               (tg2_1_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_2_1_rresp               (tg2_1_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_2_1_rlast               (tg2_1_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_2_1_rvalid              (tg2_1_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_2_1_rready              (tg2_1_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_3_0_awid                (tg3_0_axi_awid),                                   //   input,    width = 7,             axi_3_0.awid
		.axi_3_0_awaddr              (tg3_0_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_3_0_awlen               (tg3_0_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_3_0_awsize              (tg3_0_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_3_0_awburst             (tg3_0_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_3_0_awprot              (tg3_0_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_3_0_awqos               (tg3_0_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_3_0_awuser              (tg3_0_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_3_0_awvalid             (tg3_0_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_3_0_awready             (tg3_0_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_3_0_wdata               (tg3_0_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_3_0_wstrb               (tg3_0_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_3_0_wlast               (tg3_0_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_3_0_wvalid              (tg3_0_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_3_0_wready              (tg3_0_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_3_0_bid                 (tg3_0_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_3_0_bresp               (tg3_0_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_3_0_bvalid              (tg3_0_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_3_0_bready              (tg3_0_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_3_0_arid                (tg3_0_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_3_0_araddr              (tg3_0_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_3_0_arlen               (tg3_0_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_3_0_arsize              (tg3_0_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_3_0_arburst             (tg3_0_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_3_0_arprot              (tg3_0_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_3_0_arqos               (tg3_0_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_3_0_aruser              (tg3_0_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_3_0_arvalid             (tg3_0_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_3_0_arready             (tg3_0_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_3_0_rid                 (tg3_0_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_3_0_rdata               (tg3_0_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_3_0_rresp               (tg3_0_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_3_0_rlast               (tg3_0_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_3_0_rvalid              (tg3_0_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_3_0_rready              (tg3_0_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_3_1_awid                (tg3_1_axi_awid),                                   //   input,    width = 7,             axi_3_1.awid
		.axi_3_1_awaddr              (tg3_1_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_3_1_awlen               (tg3_1_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_3_1_awsize              (tg3_1_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_3_1_awburst             (tg3_1_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_3_1_awprot              (tg3_1_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_3_1_awqos               (tg3_1_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_3_1_awuser              (tg3_1_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_3_1_awvalid             (tg3_1_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_3_1_awready             (tg3_1_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_3_1_wdata               (tg3_1_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_3_1_wstrb               (tg3_1_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_3_1_wlast               (tg3_1_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_3_1_wvalid              (tg3_1_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_3_1_wready              (tg3_1_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_3_1_bid                 (tg3_1_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_3_1_bresp               (tg3_1_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_3_1_bvalid              (tg3_1_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_3_1_bready              (tg3_1_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_3_1_arid                (tg3_1_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_3_1_araddr              (tg3_1_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_3_1_arlen               (tg3_1_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_3_1_arsize              (tg3_1_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_3_1_arburst             (tg3_1_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_3_1_arprot              (tg3_1_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_3_1_arqos               (tg3_1_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_3_1_aruser              (tg3_1_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_3_1_arvalid             (tg3_1_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_3_1_arready             (tg3_1_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_3_1_rid                 (tg3_1_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_3_1_rdata               (tg3_1_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_3_1_rresp               (tg3_1_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_3_1_rlast               (tg3_1_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_3_1_rvalid              (tg3_1_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_3_1_rready              (tg3_1_axi_rready),                                 //   input,    width = 1,                    .rready
		.wmc_clk_2                   (hbm_0_example_design_wmc_clk_2_clk),               //  output,    width = 1,           wmc_clk_2.clk
		.wmcrst_n_2                  (hbm_0_example_design_wmcrst_n_2_reset),            //  output,    width = 1,          wmcrst_n_2.reset_n
		.phy_clk_4_clk               (),                                                 //  output,    width = 1,           phy_clk_4.clk
		.axi_extra_4_0_ruser_err_dbe (hbm_0_example_design_axi_extra_4_0_ruser_err_dbe), //  output,    width = 1,       axi_extra_4_0.ruser_err_dbe
		.axi_extra_4_0_ruser_data    (hbm_0_example_design_axi_extra_4_0_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_4_0_wuser_data    (tg4_0_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_4_0_wuser_strb    (tg4_0_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_4_1_ruser_err_dbe (hbm_0_example_design_axi_extra_4_1_ruser_err_dbe), //  output,    width = 1,       axi_extra_4_1.ruser_err_dbe
		.axi_extra_4_1_ruser_data    (hbm_0_example_design_axi_extra_4_1_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_4_1_wuser_data    (tg4_1_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_4_1_wuser_strb    (tg4_1_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_5_0_ruser_err_dbe (hbm_0_example_design_axi_extra_5_0_ruser_err_dbe), //  output,    width = 1,       axi_extra_5_0.ruser_err_dbe
		.axi_extra_5_0_ruser_data    (hbm_0_example_design_axi_extra_5_0_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_5_0_wuser_data    (tg5_0_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_5_0_wuser_strb    (tg5_0_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_5_1_ruser_err_dbe (hbm_0_example_design_axi_extra_5_1_ruser_err_dbe), //  output,    width = 1,       axi_extra_5_1.ruser_err_dbe
		.axi_extra_5_1_ruser_data    (hbm_0_example_design_axi_extra_5_1_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_5_1_wuser_data    (tg5_1_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_5_1_wuser_strb    (tg5_1_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.apb_4_ur_paddr              (tg4_0_apb_ur_paddr),                               //   input,   width = 16,               apb_4.ur_paddr
		.apb_4_ur_psel               (tg4_0_apb_ur_psel),                                //   input,    width = 1,                    .ur_psel
		.apb_4_ur_penable            (tg4_0_apb_ur_penable),                             //   input,    width = 1,                    .ur_penable
		.apb_4_ur_pwrite             (tg4_0_apb_ur_pwrite),                              //   input,    width = 1,                    .ur_pwrite
		.apb_4_ur_pwdata             (tg4_0_apb_ur_pwdata),                              //   input,   width = 16,                    .ur_pwdata
		.apb_4_ur_pstrb              (tg4_0_apb_ur_pstrb),                               //   input,    width = 2,                    .ur_pstrb
		.apb_4_ur_prready            (hbm_0_example_design_apb_4_ur_prready),            //  output,    width = 1,                    .ur_prready
		.apb_4_ur_prdata             (hbm_0_example_design_apb_4_ur_prdata),             //  output,   width = 16,                    .ur_prdata
		.apb_5_ur_paddr              (tg5_0_apb_ur_paddr),                               //   input,   width = 16,               apb_5.ur_paddr
		.apb_5_ur_psel               (tg5_0_apb_ur_psel),                                //   input,    width = 1,                    .ur_psel
		.apb_5_ur_penable            (tg5_0_apb_ur_penable),                             //   input,    width = 1,                    .ur_penable
		.apb_5_ur_pwrite             (tg5_0_apb_ur_pwrite),                              //   input,    width = 1,                    .ur_pwrite
		.apb_5_ur_pwdata             (tg5_0_apb_ur_pwdata),                              //   input,   width = 16,                    .ur_pwdata
		.apb_5_ur_pstrb              (tg5_0_apb_ur_pstrb),                               //   input,    width = 2,                    .ur_pstrb
		.apb_5_ur_prready            (hbm_0_example_design_apb_5_ur_prready),            //  output,    width = 1,                    .ur_prready
		.apb_5_ur_prdata             (hbm_0_example_design_apb_5_ur_prdata),             //  output,   width = 16,                    .ur_prdata
		.axi_4_0_awid                (tg4_0_axi_awid),                                   //   input,    width = 7,             axi_4_0.awid
		.axi_4_0_awaddr              (tg4_0_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_4_0_awlen               (tg4_0_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_4_0_awsize              (tg4_0_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_4_0_awburst             (tg4_0_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_4_0_awprot              (tg4_0_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_4_0_awqos               (tg4_0_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_4_0_awuser              (tg4_0_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_4_0_awvalid             (tg4_0_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_4_0_awready             (tg4_0_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_4_0_wdata               (tg4_0_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_4_0_wstrb               (tg4_0_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_4_0_wlast               (tg4_0_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_4_0_wvalid              (tg4_0_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_4_0_wready              (tg4_0_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_4_0_bid                 (tg4_0_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_4_0_bresp               (tg4_0_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_4_0_bvalid              (tg4_0_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_4_0_bready              (tg4_0_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_4_0_arid                (tg4_0_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_4_0_araddr              (tg4_0_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_4_0_arlen               (tg4_0_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_4_0_arsize              (tg4_0_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_4_0_arburst             (tg4_0_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_4_0_arprot              (tg4_0_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_4_0_arqos               (tg4_0_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_4_0_aruser              (tg4_0_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_4_0_arvalid             (tg4_0_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_4_0_arready             (tg4_0_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_4_0_rid                 (tg4_0_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_4_0_rdata               (tg4_0_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_4_0_rresp               (tg4_0_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_4_0_rlast               (tg4_0_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_4_0_rvalid              (tg4_0_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_4_0_rready              (tg4_0_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_4_1_awid                (tg4_1_axi_awid),                                   //   input,    width = 7,             axi_4_1.awid
		.axi_4_1_awaddr              (tg4_1_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_4_1_awlen               (tg4_1_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_4_1_awsize              (tg4_1_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_4_1_awburst             (tg4_1_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_4_1_awprot              (tg4_1_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_4_1_awqos               (tg4_1_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_4_1_awuser              (tg4_1_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_4_1_awvalid             (tg4_1_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_4_1_awready             (tg4_1_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_4_1_wdata               (tg4_1_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_4_1_wstrb               (tg4_1_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_4_1_wlast               (tg4_1_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_4_1_wvalid              (tg4_1_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_4_1_wready              (tg4_1_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_4_1_bid                 (tg4_1_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_4_1_bresp               (tg4_1_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_4_1_bvalid              (tg4_1_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_4_1_bready              (tg4_1_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_4_1_arid                (tg4_1_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_4_1_araddr              (tg4_1_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_4_1_arlen               (tg4_1_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_4_1_arsize              (tg4_1_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_4_1_arburst             (tg4_1_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_4_1_arprot              (tg4_1_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_4_1_arqos               (tg4_1_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_4_1_aruser              (tg4_1_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_4_1_arvalid             (tg4_1_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_4_1_arready             (tg4_1_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_4_1_rid                 (tg4_1_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_4_1_rdata               (tg4_1_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_4_1_rresp               (tg4_1_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_4_1_rlast               (tg4_1_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_4_1_rvalid              (tg4_1_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_4_1_rready              (tg4_1_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_5_0_awid                (tg5_0_axi_awid),                                   //   input,    width = 7,             axi_5_0.awid
		.axi_5_0_awaddr              (tg5_0_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_5_0_awlen               (tg5_0_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_5_0_awsize              (tg5_0_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_5_0_awburst             (tg5_0_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_5_0_awprot              (tg5_0_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_5_0_awqos               (tg5_0_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_5_0_awuser              (tg5_0_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_5_0_awvalid             (tg5_0_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_5_0_awready             (tg5_0_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_5_0_wdata               (tg5_0_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_5_0_wstrb               (tg5_0_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_5_0_wlast               (tg5_0_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_5_0_wvalid              (tg5_0_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_5_0_wready              (tg5_0_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_5_0_bid                 (tg5_0_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_5_0_bresp               (tg5_0_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_5_0_bvalid              (tg5_0_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_5_0_bready              (tg5_0_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_5_0_arid                (tg5_0_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_5_0_araddr              (tg5_0_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_5_0_arlen               (tg5_0_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_5_0_arsize              (tg5_0_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_5_0_arburst             (tg5_0_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_5_0_arprot              (tg5_0_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_5_0_arqos               (tg5_0_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_5_0_aruser              (tg5_0_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_5_0_arvalid             (tg5_0_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_5_0_arready             (tg5_0_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_5_0_rid                 (tg5_0_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_5_0_rdata               (tg5_0_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_5_0_rresp               (tg5_0_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_5_0_rlast               (tg5_0_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_5_0_rvalid              (tg5_0_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_5_0_rready              (tg5_0_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_5_1_awid                (tg5_1_axi_awid),                                   //   input,    width = 7,             axi_5_1.awid
		.axi_5_1_awaddr              (tg5_1_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_5_1_awlen               (tg5_1_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_5_1_awsize              (tg5_1_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_5_1_awburst             (tg5_1_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_5_1_awprot              (tg5_1_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_5_1_awqos               (tg5_1_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_5_1_awuser              (tg5_1_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_5_1_awvalid             (tg5_1_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_5_1_awready             (tg5_1_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_5_1_wdata               (tg5_1_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_5_1_wstrb               (tg5_1_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_5_1_wlast               (tg5_1_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_5_1_wvalid              (tg5_1_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_5_1_wready              (tg5_1_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_5_1_bid                 (tg5_1_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_5_1_bresp               (tg5_1_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_5_1_bvalid              (tg5_1_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_5_1_bready              (tg5_1_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_5_1_arid                (tg5_1_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_5_1_araddr              (tg5_1_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_5_1_arlen               (tg5_1_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_5_1_arsize              (tg5_1_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_5_1_arburst             (tg5_1_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_5_1_arprot              (tg5_1_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_5_1_arqos               (tg5_1_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_5_1_aruser              (tg5_1_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_5_1_arvalid             (tg5_1_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_5_1_arready             (tg5_1_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_5_1_rid                 (tg5_1_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_5_1_rdata               (tg5_1_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_5_1_rresp               (tg5_1_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_5_1_rlast               (tg5_1_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_5_1_rvalid              (tg5_1_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_5_1_rready              (tg5_1_axi_rready),                                 //   input,    width = 1,                    .rready
		.wmc_clk_4                   (hbm_0_example_design_wmc_clk_4_clk),               //  output,    width = 1,           wmc_clk_4.clk
		.wmcrst_n_4                  (hbm_0_example_design_wmcrst_n_4_reset),            //  output,    width = 1,          wmcrst_n_4.reset_n
		.phy_clk_6_clk               (),                                                 //  output,    width = 1,           phy_clk_6.clk
		.axi_extra_6_0_ruser_err_dbe (hbm_0_example_design_axi_extra_6_0_ruser_err_dbe), //  output,    width = 1,       axi_extra_6_0.ruser_err_dbe
		.axi_extra_6_0_ruser_data    (hbm_0_example_design_axi_extra_6_0_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_6_0_wuser_data    (tg6_0_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_6_0_wuser_strb    (tg6_0_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_6_1_ruser_err_dbe (hbm_0_example_design_axi_extra_6_1_ruser_err_dbe), //  output,    width = 1,       axi_extra_6_1.ruser_err_dbe
		.axi_extra_6_1_ruser_data    (hbm_0_example_design_axi_extra_6_1_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_6_1_wuser_data    (tg6_1_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_6_1_wuser_strb    (tg6_1_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_7_0_ruser_err_dbe (hbm_0_example_design_axi_extra_7_0_ruser_err_dbe), //  output,    width = 1,       axi_extra_7_0.ruser_err_dbe
		.axi_extra_7_0_ruser_data    (hbm_0_example_design_axi_extra_7_0_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_7_0_wuser_data    (tg7_0_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_7_0_wuser_strb    (tg7_0_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.axi_extra_7_1_ruser_err_dbe (hbm_0_example_design_axi_extra_7_1_ruser_err_dbe), //  output,    width = 1,       axi_extra_7_1.ruser_err_dbe
		.axi_extra_7_1_ruser_data    (hbm_0_example_design_axi_extra_7_1_ruser_data),    //  output,   width = 32,                    .ruser_data
		.axi_extra_7_1_wuser_data    (tg7_1_axi_extra_wuser_data),                       //   input,   width = 32,                    .wuser_data
		.axi_extra_7_1_wuser_strb    (tg7_1_axi_extra_wuser_strb),                       //   input,    width = 4,                    .wuser_strb
		.apb_6_ur_paddr              (tg6_0_apb_ur_paddr),                               //   input,   width = 16,               apb_6.ur_paddr
		.apb_6_ur_psel               (tg6_0_apb_ur_psel),                                //   input,    width = 1,                    .ur_psel
		.apb_6_ur_penable            (tg6_0_apb_ur_penable),                             //   input,    width = 1,                    .ur_penable
		.apb_6_ur_pwrite             (tg6_0_apb_ur_pwrite),                              //   input,    width = 1,                    .ur_pwrite
		.apb_6_ur_pwdata             (tg6_0_apb_ur_pwdata),                              //   input,   width = 16,                    .ur_pwdata
		.apb_6_ur_pstrb              (tg6_0_apb_ur_pstrb),                               //   input,    width = 2,                    .ur_pstrb
		.apb_6_ur_prready            (hbm_0_example_design_apb_6_ur_prready),            //  output,    width = 1,                    .ur_prready
		.apb_6_ur_prdata             (hbm_0_example_design_apb_6_ur_prdata),             //  output,   width = 16,                    .ur_prdata
		.apb_7_ur_paddr              (tg7_0_apb_ur_paddr),                               //   input,   width = 16,               apb_7.ur_paddr
		.apb_7_ur_psel               (tg7_0_apb_ur_psel),                                //   input,    width = 1,                    .ur_psel
		.apb_7_ur_penable            (tg7_0_apb_ur_penable),                             //   input,    width = 1,                    .ur_penable
		.apb_7_ur_pwrite             (tg7_0_apb_ur_pwrite),                              //   input,    width = 1,                    .ur_pwrite
		.apb_7_ur_pwdata             (tg7_0_apb_ur_pwdata),                              //   input,   width = 16,                    .ur_pwdata
		.apb_7_ur_pstrb              (tg7_0_apb_ur_pstrb),                               //   input,    width = 2,                    .ur_pstrb
		.apb_7_ur_prready            (hbm_0_example_design_apb_7_ur_prready),            //  output,    width = 1,                    .ur_prready
		.apb_7_ur_prdata             (hbm_0_example_design_apb_7_ur_prdata),             //  output,   width = 16,                    .ur_prdata
		.axi_6_0_awid                (tg6_0_axi_awid),                                   //   input,    width = 7,             axi_6_0.awid
		.axi_6_0_awaddr              (tg6_0_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_6_0_awlen               (tg6_0_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_6_0_awsize              (tg6_0_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_6_0_awburst             (tg6_0_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_6_0_awprot              (tg6_0_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_6_0_awqos               (tg6_0_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_6_0_awuser              (tg6_0_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_6_0_awvalid             (tg6_0_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_6_0_awready             (tg6_0_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_6_0_wdata               (tg6_0_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_6_0_wstrb               (tg6_0_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_6_0_wlast               (tg6_0_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_6_0_wvalid              (tg6_0_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_6_0_wready              (tg6_0_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_6_0_bid                 (tg6_0_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_6_0_bresp               (tg6_0_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_6_0_bvalid              (tg6_0_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_6_0_bready              (tg6_0_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_6_0_arid                (tg6_0_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_6_0_araddr              (tg6_0_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_6_0_arlen               (tg6_0_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_6_0_arsize              (tg6_0_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_6_0_arburst             (tg6_0_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_6_0_arprot              (tg6_0_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_6_0_arqos               (tg6_0_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_6_0_aruser              (tg6_0_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_6_0_arvalid             (tg6_0_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_6_0_arready             (tg6_0_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_6_0_rid                 (tg6_0_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_6_0_rdata               (tg6_0_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_6_0_rresp               (tg6_0_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_6_0_rlast               (tg6_0_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_6_0_rvalid              (tg6_0_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_6_0_rready              (tg6_0_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_6_1_awid                (tg6_1_axi_awid),                                   //   input,    width = 7,             axi_6_1.awid
		.axi_6_1_awaddr              (tg6_1_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_6_1_awlen               (tg6_1_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_6_1_awsize              (tg6_1_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_6_1_awburst             (tg6_1_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_6_1_awprot              (tg6_1_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_6_1_awqos               (tg6_1_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_6_1_awuser              (tg6_1_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_6_1_awvalid             (tg6_1_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_6_1_awready             (tg6_1_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_6_1_wdata               (tg6_1_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_6_1_wstrb               (tg6_1_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_6_1_wlast               (tg6_1_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_6_1_wvalid              (tg6_1_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_6_1_wready              (tg6_1_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_6_1_bid                 (tg6_1_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_6_1_bresp               (tg6_1_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_6_1_bvalid              (tg6_1_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_6_1_bready              (tg6_1_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_6_1_arid                (tg6_1_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_6_1_araddr              (tg6_1_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_6_1_arlen               (tg6_1_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_6_1_arsize              (tg6_1_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_6_1_arburst             (tg6_1_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_6_1_arprot              (tg6_1_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_6_1_arqos               (tg6_1_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_6_1_aruser              (tg6_1_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_6_1_arvalid             (tg6_1_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_6_1_arready             (tg6_1_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_6_1_rid                 (tg6_1_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_6_1_rdata               (tg6_1_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_6_1_rresp               (tg6_1_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_6_1_rlast               (tg6_1_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_6_1_rvalid              (tg6_1_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_6_1_rready              (tg6_1_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_7_0_awid                (tg7_0_axi_awid),                                   //   input,    width = 7,             axi_7_0.awid
		.axi_7_0_awaddr              (tg7_0_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_7_0_awlen               (tg7_0_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_7_0_awsize              (tg7_0_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_7_0_awburst             (tg7_0_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_7_0_awprot              (tg7_0_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_7_0_awqos               (tg7_0_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_7_0_awuser              (tg7_0_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_7_0_awvalid             (tg7_0_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_7_0_awready             (tg7_0_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_7_0_wdata               (tg7_0_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_7_0_wstrb               (tg7_0_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_7_0_wlast               (tg7_0_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_7_0_wvalid              (tg7_0_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_7_0_wready              (tg7_0_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_7_0_bid                 (tg7_0_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_7_0_bresp               (tg7_0_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_7_0_bvalid              (tg7_0_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_7_0_bready              (tg7_0_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_7_0_arid                (tg7_0_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_7_0_araddr              (tg7_0_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_7_0_arlen               (tg7_0_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_7_0_arsize              (tg7_0_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_7_0_arburst             (tg7_0_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_7_0_arprot              (tg7_0_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_7_0_arqos               (tg7_0_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_7_0_aruser              (tg7_0_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_7_0_arvalid             (tg7_0_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_7_0_arready             (tg7_0_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_7_0_rid                 (tg7_0_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_7_0_rdata               (tg7_0_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_7_0_rresp               (tg7_0_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_7_0_rlast               (tg7_0_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_7_0_rvalid              (tg7_0_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_7_0_rready              (tg7_0_axi_rready),                                 //   input,    width = 1,                    .rready
		.axi_7_1_awid                (tg7_1_axi_awid),                                   //   input,    width = 7,             axi_7_1.awid
		.axi_7_1_awaddr              (tg7_1_axi_awaddr),                                 //   input,   width = 30,                    .awaddr
		.axi_7_1_awlen               (tg7_1_axi_awlen),                                  //   input,    width = 8,                    .awlen
		.axi_7_1_awsize              (tg7_1_axi_awsize),                                 //   input,    width = 3,                    .awsize
		.axi_7_1_awburst             (tg7_1_axi_awburst),                                //   input,    width = 2,                    .awburst
		.axi_7_1_awprot              (tg7_1_axi_awprot),                                 //   input,    width = 3,                    .awprot
		.axi_7_1_awqos               (tg7_1_axi_awqos),                                  //   input,    width = 4,                    .awqos
		.axi_7_1_awuser              (tg7_1_axi_awuser),                                 //   input,    width = 1,                    .awuser
		.axi_7_1_awvalid             (tg7_1_axi_awvalid),                                //   input,    width = 1,                    .awvalid
		.axi_7_1_awready             (tg7_1_axi_awready),                                //  output,    width = 1,                    .awready
		.axi_7_1_wdata               (tg7_1_axi_wdata),                                  //   input,  width = 256,                    .wdata
		.axi_7_1_wstrb               (tg7_1_axi_wstrb),                                  //   input,   width = 32,                    .wstrb
		.axi_7_1_wlast               (tg7_1_axi_wlast),                                  //   input,    width = 1,                    .wlast
		.axi_7_1_wvalid              (tg7_1_axi_wvalid),                                 //   input,    width = 1,                    .wvalid
		.axi_7_1_wready              (tg7_1_axi_wready),                                 //  output,    width = 1,                    .wready
		.axi_7_1_bid                 (tg7_1_axi_bid),                                    //  output,    width = 7,                    .bid
		.axi_7_1_bresp               (tg7_1_axi_bresp),                                  //  output,    width = 2,                    .bresp
		.axi_7_1_bvalid              (tg7_1_axi_bvalid),                                 //  output,    width = 1,                    .bvalid
		.axi_7_1_bready              (tg7_1_axi_bready),                                 //   input,    width = 1,                    .bready
		.axi_7_1_arid                (tg7_1_axi_arid),                                   //   input,    width = 7,                    .arid
		.axi_7_1_araddr              (tg7_1_axi_araddr),                                 //   input,   width = 30,                    .araddr
		.axi_7_1_arlen               (tg7_1_axi_arlen),                                  //   input,    width = 8,                    .arlen
		.axi_7_1_arsize              (tg7_1_axi_arsize),                                 //   input,    width = 3,                    .arsize
		.axi_7_1_arburst             (tg7_1_axi_arburst),                                //   input,    width = 2,                    .arburst
		.axi_7_1_arprot              (tg7_1_axi_arprot),                                 //   input,    width = 3,                    .arprot
		.axi_7_1_arqos               (tg7_1_axi_arqos),                                  //   input,    width = 4,                    .arqos
		.axi_7_1_aruser              (tg7_1_axi_aruser),                                 //   input,    width = 1,                    .aruser
		.axi_7_1_arvalid             (tg7_1_axi_arvalid),                                //   input,    width = 1,                    .arvalid
		.axi_7_1_arready             (tg7_1_axi_arready),                                //  output,    width = 1,                    .arready
		.axi_7_1_rid                 (tg7_1_axi_rid),                                    //  output,    width = 7,                    .rid
		.axi_7_1_rdata               (tg7_1_axi_rdata),                                  //  output,  width = 256,                    .rdata
		.axi_7_1_rresp               (tg7_1_axi_rresp),                                  //  output,    width = 2,                    .rresp
		.axi_7_1_rlast               (tg7_1_axi_rlast),                                  //  output,    width = 1,                    .rlast
		.axi_7_1_rvalid              (tg7_1_axi_rvalid),                                 //  output,    width = 1,                    .rvalid
		.axi_7_1_rready              (tg7_1_axi_rready),                                 //   input,    width = 1,                    .rready
		.wmc_clk_6                   (hbm_0_example_design_wmc_clk_6_clk),               //  output,    width = 1,           wmc_clk_6.clk
		.wmcrst_n_6                  (hbm_0_example_design_wmcrst_n_6_reset)             //  output,    width = 1,          wmcrst_n_6.reset_n
	);

	ed_synth_ninit_done_splitter ninit_done_splitter (
		.sig_input     (reset_release_ip_ninit_done_ninit_done),          //   input,  width = 1,     sig_input_if.ninit_done
		.sig_output_0  (ninit_done_splitter_sig_output_if_0_ninit_done),  //  output,  width = 1,  sig_output_if_0.ninit_done
		.sig_output_1  (ninit_done_splitter_sig_output_if_1_ninit_done),  //  output,  width = 1,  sig_output_if_1.ninit_done
		.sig_output_2  (ninit_done_splitter_sig_output_if_2_ninit_done),  //  output,  width = 1,  sig_output_if_2.ninit_done
		.sig_output_3  (ninit_done_splitter_sig_output_if_3_ninit_done),  //  output,  width = 1,  sig_output_if_3.ninit_done
		.sig_output_4  (ninit_done_splitter_sig_output_if_4_ninit_done),  //  output,  width = 1,  sig_output_if_4.ninit_done
		.sig_output_5  (ninit_done_splitter_sig_output_if_5_ninit_done),  //  output,  width = 1,  sig_output_if_5.ninit_done
		.sig_output_6  (ninit_done_splitter_sig_output_if_6_ninit_done),  //  output,  width = 1,  sig_output_if_6.ninit_done
		.sig_output_7  (ninit_done_splitter_sig_output_if_7_ninit_done),  //  output,  width = 1,  sig_output_if_7.ninit_done
		.sig_output_8  (ninit_done_splitter_sig_output_if_8_ninit_done),  //  output,  width = 1,  sig_output_if_8.ninit_done
		.sig_output_9  (ninit_done_splitter_sig_output_if_9_ninit_done),  //  output,  width = 1,  sig_output_if_9.ninit_done
		.sig_output_10 (ninit_done_splitter_sig_output_if_10_ninit_done), //  output,  width = 1, sig_output_if_10.ninit_done
		.sig_output_11 (ninit_done_splitter_sig_output_if_11_ninit_done), //  output,  width = 1, sig_output_if_11.ninit_done
		.sig_output_12 (ninit_done_splitter_sig_output_if_12_ninit_done), //  output,  width = 1, sig_output_if_12.ninit_done
		.sig_output_13 (ninit_done_splitter_sig_output_if_13_ninit_done), //  output,  width = 1, sig_output_if_13.ninit_done
		.sig_output_14 (ninit_done_splitter_sig_output_if_14_ninit_done), //  output,  width = 1, sig_output_if_14.ninit_done
		.sig_output_15 (ninit_done_splitter_sig_output_if_15_ninit_done)  //  output,  width = 1, sig_output_if_15.ninit_done
	);

	ed_synth_reset_release_ip reset_release_ip (
		.ninit_done (reset_release_ip_ninit_done_ninit_done)  //  output,  width = 1, ninit_done.ninit_done
	);

	assign tg0_0_apb_ur_paddr = 0;
	assign tg0_0_apb_ur_psel = 0;
	assign tg0_0_apb_ur_penable = 0;
	assign tg0_0_apb_ur_pwrite = 0;
	assign tg0_0_apb_ur_pwdata = 0;
	assign tg0_0_apb_ur_pstrb = 0;
	assign tg0_1_apb_ur_paddr = 0;
	assign tg0_1_apb_ur_psel = 0;
	assign tg0_1_apb_ur_penable = 0;
	assign tg0_1_apb_ur_pwrite = 0;
	assign tg0_1_apb_ur_pwdata = 0;
	assign tg0_1_apb_ur_pstrb = 0;
	assign tg1_0_apb_ur_paddr = 0;
	assign tg1_0_apb_ur_psel = 0;
	assign tg1_0_apb_ur_penable = 0;
	assign tg1_0_apb_ur_pwrite = 0;
	assign tg1_0_apb_ur_pwdata = 0;
	assign tg1_0_apb_ur_pstrb = 0;
	assign tg1_1_apb_ur_paddr = 0;
	assign tg1_1_apb_ur_psel = 0;
	assign tg1_1_apb_ur_penable = 0;
	assign tg1_1_apb_ur_pwrite = 0;
	assign tg1_1_apb_ur_pwdata = 0;
	assign tg1_1_apb_ur_pstrb = 0;
	assign tg2_0_apb_ur_paddr = 0;
	assign tg2_0_apb_ur_psel = 0;
	assign tg2_0_apb_ur_penable = 0;
	assign tg2_0_apb_ur_pwrite = 0;
	assign tg2_0_apb_ur_pwdata = 0;
	assign tg2_0_apb_ur_pstrb = 0;
	assign tg2_1_apb_ur_paddr = 0;
	assign tg2_1_apb_ur_psel = 0;
	assign tg2_1_apb_ur_penable = 0;
	assign tg2_1_apb_ur_pwrite = 0;
	assign tg2_1_apb_ur_pwdata = 0;
	assign tg2_1_apb_ur_pstrb = 0;
	assign tg3_0_apb_ur_paddr = 0;
	assign tg3_0_apb_ur_psel = 0;
	assign tg3_0_apb_ur_penable = 0;
	assign tg3_0_apb_ur_pwrite = 0;
	assign tg3_0_apb_ur_pwdata = 0;
	assign tg3_0_apb_ur_pstrb = 0;
	assign tg3_1_apb_ur_paddr = 0;
	assign tg3_1_apb_ur_psel = 0;
	assign tg3_1_apb_ur_penable = 0;
	assign tg3_1_apb_ur_pwrite = 0;
	assign tg3_1_apb_ur_pwdata = 0;
	assign tg3_1_apb_ur_pstrb = 0;
	assign tg4_0_apb_ur_paddr = 0;
	assign tg4_0_apb_ur_psel = 0;
	assign tg4_0_apb_ur_penable = 0;
	assign tg4_0_apb_ur_pwrite = 0;
	assign tg4_0_apb_ur_pwdata = 0;
	assign tg4_0_apb_ur_pstrb = 0;
	assign tg4_1_apb_ur_paddr = 0;
	assign tg4_1_apb_ur_psel = 0;
	assign tg4_1_apb_ur_penable = 0;
	assign tg4_1_apb_ur_pwrite = 0;
	assign tg4_1_apb_ur_pwdata = 0;
	assign tg4_1_apb_ur_pstrb = 0;
	assign tg5_0_apb_ur_paddr = 0;
	assign tg5_0_apb_ur_psel = 0;
	assign tg5_0_apb_ur_penable = 0;
	assign tg5_0_apb_ur_pwrite = 0;
	assign tg5_0_apb_ur_pwdata = 0;
	assign tg5_0_apb_ur_pstrb = 0;
	assign tg5_1_apb_ur_paddr = 0;
	assign tg5_1_apb_ur_psel = 0;
	assign tg5_1_apb_ur_penable = 0;
	assign tg5_1_apb_ur_pwrite = 0;
	assign tg5_1_apb_ur_pwdata = 0;
	assign tg5_1_apb_ur_pstrb = 0;
	assign tg6_0_apb_ur_paddr = 0;
	assign tg6_0_apb_ur_psel = 0;
	assign tg6_0_apb_ur_penable = 0;
	assign tg6_0_apb_ur_pwrite = 0;
	assign tg6_0_apb_ur_pwdata = 0;
	assign tg6_0_apb_ur_pstrb = 0;
	assign tg6_1_apb_ur_paddr = 0;
	assign tg6_1_apb_ur_psel = 0;
	assign tg6_1_apb_ur_penable = 0;
	assign tg6_1_apb_ur_pwrite = 0;
	assign tg6_1_apb_ur_pwdata = 0;
	assign tg6_1_apb_ur_pstrb = 0;
	assign tg7_0_apb_ur_paddr = 0;
	assign tg7_0_apb_ur_psel = 0;
	assign tg7_0_apb_ur_penable = 0;
	assign tg7_0_apb_ur_pwrite = 0;
	assign tg7_0_apb_ur_pwdata = 0;
	assign tg7_0_apb_ur_pstrb = 0;
	assign tg7_1_apb_ur_paddr = 0;
	assign tg7_1_apb_ur_psel = 0;
	assign tg7_1_apb_ur_penable = 0;
	assign tg7_1_apb_ur_pwrite = 0;
	assign tg7_1_apb_ur_pwdata = 0;
	assign tg7_1_apb_ur_pstrb = 0;

  FGPU uut(
    .clk(hbm_0_example_design_wmc_clk_0_clk),
    //slave axi {{{
    .s0_awaddr(s0_awaddr),
    .s0_awprot(s0_awprot),
    .s0_awvalid(s0_awvalid),
    .s0_awready(s0_awready),
  
    .s0_wdata(s0_wdata),
    .s0_wstrb(s0_wstrb),
    .s0_wvalid(s0_wvalid),
    .s0_wready(s0_wready),
  
    .s0_bresp(s0_bresp),
    .s0_bvalid(s0_bvalid),
    .s0_bready(s0_bready),
  
    .s0_araddr(s0_araddr),
    .s0_arprot(s0_arprot),
    .s0_arvalid(s0_arvalid),
    .s0_arready(s0_arready),
  
    .s0_rdata(s0_rdata),
    .s0_rresp(s0_rresp),
    .s0_rvalid(s0_rvalid),
    .s0_rready(s0_rready),
    //-- }}}
    //-- axi master 0 {{{
    //-- ar channel
    .m0_araddr(m0_araddr),
    .m0_arlen(m0_arlen),
    .m0_arsize(m0_arsize),
    .m0_arburst(m0_arburst),
    .m0_arvalid(m0_arvalid),
    .m0_arready(m0_arready),
    .m0_arid(m0_arid),
    //-- r channel
    .m0_rdata(m0_rdata),
    .m0_rresp(m0_rresp),
    .m0_rlast(m0_rlast),
    .m0_rvalid(m0_rvalid),
    .m0_rready(m0_rready),
    .m0_rid(m0_rid),
    //-- aw channel
    .m0_awvalid(m0_awvalid),
    .m0_awaddr(m0_awaddr),
    .m0_awready(m0_awready),
    .m0_awlen(m0_awlen),
    .m0_awsize(m0_awsize),
    .m0_awburst(m0_awburst),
    .m0_awid(m0_awid),
    //--    .w channel
    .m0_wdata(m0_wdata),
    .m0_wstrb(m0_wstrb),
    .m0_wlast(m0_wlast),
    .m0_wvalid(m0_wvalid),
    .m0_wready(m0_wready),
    //-- bchannel
    .m0_bvalid(m0_bvalid),
    .m0_bready(m0_bready),
    .m0_bid(m0_bid),
    //-- }}}
    //-- interface 1 {{{
    //-- ar channel
    .m1_araddr(m1_araddr),
    .m1_arlen(m1_arlen),
    .m1_arsize(m1_arsize),
    .m1_arburst(m1_arburst),
    .m1_arvalid(m1_arvalid),
    .m1_arready(m1_arready),
    .m1_arid(m1_arid),
    //-- r channel
    .m1_rdata(m1_rdata),
    .m1_rresp(m1_rresp),
    .m1_rlast(m1_rlast),
    .m1_rvalid(m1_rvalid),
    .m1_rready(m1_rready),
    .m1_rid(m1_rid),
    //-- aw channel
    .m1_awvalid(m1_awvalid),
    .m1_awaddr(m1_awaddr),
    .m1_awready(m1_awready),
    .m1_awlen(m1_awlen),
    .m1_awsize(m1_awsize),
    .m1_awburst(m1_awburst),
    .m1_awid(m1_awid),
    //-- w channel
    .m1_wdata(m1_wdata),
    .m1_wstrb(m1_wstrb),
    .m1_wlast(m1_wlast),
    .m1_wvalid(m1_wvalid),
    .m1_wready(m1_wready),
    //-- b channel
    .m1_bready(m1_bready),
    .m1_bvalid(m1_bvalid),
    .m1_bid(m1_bid),
    //--}}}
    //-- interface 2 {{{
    //-- ar channel
    .m2_araddr(m2_araddr),
    .m2_arlen(m2_arlen),
    .m2_arsize(m2_arsize),
    .m2_arburst(m2_arburst),
    .m2_arvalid(m2_arvalid),
    .m2_arready(m2_arready),
    .m2_arid(m2_arid),
    //-- r channel
    .m2_rdata(m2_rdata),
    .m2_rresp(m2_rresp),
    .m2_rlast(m2_rlast),
    .m2_rvalid(m2_rvalid),
    .m2_rready(m2_rready),
    .m2_rid(m2_rid),
    //-- aw channel
    .m2_awvalid(m2_awvalid),
    .m2_awaddr(m2_awaddr),
    .m2_awready(m2_awready),
    .m2_awlen(m2_awlen),
    .m2_awsize(m2_awsize),
    .m2_awburst(m2_awburst),
    .m2_awid(m2_awid),
    //-- w channel
    .m2_wdata(m2_wdata),
    .m2_wstrb(m2_wstrb),
    .m2_wlast(m2_wlast),
    .m2_wvalid(m2_wvalid),
    .m2_wready(m2_wready),
    //-- b channel
    .m2_bready(m2_bready),
    .m2_bvalid(m2_bvalid),
    .m2_bid(m2_bid),
    //--}}}
    //-- interface 3 {{{
    //-- ar channel
    .m3_araddr(m3_araddr),
    .m3_arlen(m3_arlen),
    .m3_arsize(m3_arsize),
    .m3_arburst(m3_arburst),
    .m3_arvalid(m3_arvalid),
    .m3_arready(m3_arready),
    .m3_arid(m3_arid),
    //-- r channel
    .m3_rdata(m3_rdata),
    .m3_rresp(m3_rresp),
    .m3_rlast(m3_rlast),
    .m3_rvalid(m3_rvalid),
    .m3_rready(m3_rready),
    .m3_rid(m3_rid),
    //-- aw channel
    .m3_awvalid(m3_awvalid),
    .m3_awaddr(m3_awaddr),
    .m3_awready(m3_awready),
    .m3_awlen(m3_awlen),
    .m3_awsize(m3_awsize),
    .m3_awburst(m3_awburst),
    .m3_awid(m3_awid),
    //-- w channel
    .m3_wdata(m3_wdata),
    .m3_wstrb(m3_wstrb),
    .m3_wlast(m3_wlast),
    .m3_wvalid(m3_wvalid),
    .m3_wready(m3_wready),
    //-- b channel
    .m3_bready(m3_bready),
    .m3_bvalid(m3_bvalid),
    .m3_bid(m3_bid),

    .nrst(hbm_0_example_design_wmcrst_n_0_reset)
  );

  assign tg0_0_axi_rready = tg0_0_axi_rvalid & tg2_0_axi_rvalid & tg4_0_axi_rvalid & tg6_0_axi_rvalid;
  assign tg2_0_axi_rready = tg0_0_axi_rvalid & tg2_0_axi_rvalid & tg4_0_axi_rvalid & tg6_0_axi_rvalid;
  assign tg4_0_axi_rready = tg0_0_axi_rvalid & tg2_0_axi_rvalid & tg4_0_axi_rvalid & tg6_0_axi_rvalid;
  assign tg6_0_axi_rready = tg0_0_axi_rvalid & tg2_0_axi_rvalid & tg4_0_axi_rvalid & tg6_0_axi_rvalid;
  assign tg0_1_axi_rready = tg0_1_axi_rvalid & tg2_1_axi_rvalid & tg4_1_axi_rvalid & tg6_1_axi_rvalid;
  assign tg2_1_axi_rready = tg0_1_axi_rvalid & tg2_1_axi_rvalid & tg4_1_axi_rvalid & tg6_1_axi_rvalid;
  assign tg4_1_axi_rready = tg0_1_axi_rvalid & tg2_1_axi_rvalid & tg4_1_axi_rvalid & tg6_1_axi_rvalid;
  assign tg6_1_axi_rready = tg0_1_axi_rvalid & tg2_1_axi_rvalid & tg4_1_axi_rvalid & tg6_1_axi_rvalid;
  assign tg1_0_axi_rready = tg1_0_axi_rvalid & tg3_0_axi_rvalid & tg5_0_axi_rvalid & tg7_0_axi_rvalid;
  assign tg3_0_axi_rready = tg1_0_axi_rvalid & tg3_0_axi_rvalid & tg5_0_axi_rvalid & tg7_0_axi_rvalid;
  assign tg5_0_axi_rready = tg1_0_axi_rvalid & tg3_0_axi_rvalid & tg5_0_axi_rvalid & tg7_0_axi_rvalid;
  assign tg7_0_axi_rready = tg1_0_axi_rvalid & tg3_0_axi_rvalid & tg5_0_axi_rvalid & tg7_0_axi_rvalid;
  assign tg1_1_axi_rready = tg1_1_axi_rvalid & tg3_1_axi_rvalid & tg5_1_axi_rvalid & tg7_1_axi_rvalid;
  assign tg3_1_axi_rready = tg1_1_axi_rvalid & tg3_1_axi_rvalid & tg5_1_axi_rvalid & tg7_1_axi_rvalid;
  assign tg5_1_axi_rready = tg1_1_axi_rvalid & tg3_1_axi_rvalid & tg5_1_axi_rvalid & tg7_1_axi_rvalid;
  assign tg7_1_axi_rready = tg1_1_axi_rvalid & tg3_1_axi_rvalid & tg5_1_axi_rvalid & tg7_1_axi_rvalid;

  assign tg0_0_axi_awburst = m0_awburst;
  assign tg0_0_axi_awuser = 1'b0;
  assign tg0_0_axi_arlen = m0_arlen;
  assign tg0_0_axi_arqos = 4'b0;
  assign tg0_0_axi_wstrb = m0_wstrb[31:0];
  assign m0_wready = tg0_0_axi_wready & tg2_0_axi_wready & tg4_0_axi_wready & tg6_0_axi_wready;
  assign m0_rid = tg0_0_axi_rid;
  assign tg0_0_axi_awlen = m0_awlen;
  assign tg0_0_axi_awqos = 4'b0;
  assign tg0_0_axi_wvalid = m0_wvalid & m0_wready;
  assign tg0_0_axi_araddr = {m0_araddr[31:7], 5'b0};
  assign tg0_0_axi_arprot = 3'b0;
  assign tg0_0_axi_awprot = 3'b0;
  assign tg0_0_axi_wdata = m0_wdata[255:0];
  assign tg0_0_axi_arvalid = m0_arvalid & m0_arready;
  assign tg0_0_axi_arid = m0_arid;
  assign tg0_0_axi_awaddr = {m0_awaddr[31:7], 5'b0};
  assign m0_arready = tg0_0_axi_arready & tg2_0_axi_arready & tg4_0_axi_arready & tg6_0_axi_arready;
  assign m0_rdata[255:0] = tg0_0_axi_rdata;
  assign m0_awready = tg0_0_axi_awready & tg2_0_axi_awready & tg4_0_axi_awready & tg6_0_axi_awready;
  assign tg0_0_axi_arburst = m0_arburst;
  assign tg0_0_axi_arsize = m0_arsize;
  assign tg0_0_axi_bready = m0_bready;
  assign m0_rlast = tg0_0_axi_rlast;
  assign tg0_0_axi_wlast = m0_wlast;
  assign tg0_0_axi_awid = m0_awid;
  assign m0_bid = tg0_0_axi_bid;
  assign m0_bvalid = tg0_0_axi_bvalid;
  assign tg0_0_axi_awsize = m0_awsize;
  assign tg0_0_axi_awvalid = m0_awvalid & m0_awready;
  assign tg0_0_axi_aruser = 1'b0;
  assign m0_rvalid = tg0_0_axi_rvalid & tg2_0_axi_rvalid & tg4_0_axi_rvalid & tg6_0_axi_rvalid;

  assign tg2_0_axi_awburst = m0_awburst;
  assign tg2_0_axi_awuser = 1'b0;
  assign tg2_0_axi_arlen = m0_arlen;
  assign tg2_0_axi_arqos = 4'b0;
  assign tg2_0_axi_wstrb = m0_wstrb[63:32];
  assign tg2_0_axi_awlen = m0_awlen;
  assign tg2_0_axi_awqos = 4'b0;
  assign tg2_0_axi_wvalid = m0_wvalid & m0_wready;
  assign tg2_0_axi_araddr = {m0_araddr[31:7], 5'b0};
  assign tg2_0_axi_arprot = 3'b0;
  assign tg2_0_axi_awprot = 3'b0;
  assign tg2_0_axi_wdata = m0_wdata[255:0];
  assign tg2_0_axi_arvalid = m0_arvalid & m0_arready;
  assign tg2_0_axi_arid = m0_arid;
  assign tg2_0_axi_awaddr = {m0_awaddr[31:7], 5'b0};
  assign m0_rdata[511:256] = tg2_0_axi_rdata;
  assign tg2_0_axi_arburst = m0_arburst;
  assign tg2_0_axi_arsize = m0_arsize;
  assign tg2_0_axi_bready = m0_bready;
  assign tg2_0_axi_wlast = m0_wlast;
  assign tg2_0_axi_awid = m0_awid;
  assign tg2_0_axi_awsize = m0_awsize;
  assign tg2_0_axi_awvalid = m0_awvalid & m0_awready;
  assign tg2_0_axi_aruser = 1'b0;

  assign tg4_0_axi_awburst = m0_awburst;
  assign tg4_0_axi_awuser = 1'b0;
  assign tg4_0_axi_arlen = m0_arlen;
  assign tg4_0_axi_arqos = 4'b0;
  assign tg4_0_axi_wstrb = m0_wstrb[95:64];
  assign tg4_0_axi_awlen = m0_awlen;
  assign tg4_0_axi_awqos = 4'b0;
  assign tg4_0_axi_wvalid = m0_wvalid & m0_wready;
  assign tg4_0_axi_araddr = {m0_araddr[31:7], 5'b0};
  assign tg4_0_axi_arprot = 3'b0;
  assign tg4_0_axi_awprot = 3'b0;
  assign tg4_0_axi_wdata = m0_wdata[255:0];
  assign tg4_0_axi_arvalid = m0_arvalid & m0_arready;
  assign tg4_0_axi_arid = m0_arid;
  assign tg4_0_axi_awaddr = {m0_awaddr[31:7], 5'b0};
  assign m0_rdata[767:512] = tg4_0_axi_rdata;
  assign tg4_0_axi_arburst = m0_arburst;
  assign tg4_0_axi_arsize = m0_arsize;
  assign tg4_0_axi_bready = m0_bready;
  assign tg4_0_axi_wlast = m0_wlast;
  assign tg4_0_axi_awid = m0_awid;
  assign tg4_0_axi_awsize = m0_awsize;
  assign tg4_0_axi_awvalid = m0_awvalid & m0_awready;
  assign tg4_0_axi_aruser = 1'b0;

  assign tg6_0_axi_awburst = m0_awburst;
  assign tg6_0_axi_awuser = 1'b0;
  assign tg6_0_axi_arlen = m0_arlen;
  assign tg6_0_axi_arqos = 4'b0;
  assign tg6_0_axi_wstrb = m0_wstrb[127:96];
  assign tg6_0_axi_awlen = m0_awlen;
  assign tg6_0_axi_awqos = 4'b0;
  assign tg6_0_axi_wvalid = m0_wvalid & m0_wready;
  assign tg6_0_axi_araddr = {m0_araddr[31:7], 5'b0};
  assign tg6_0_axi_arprot = 3'b0;
  assign tg6_0_axi_awprot = 3'b0;
  assign tg6_0_axi_wdata = m0_wdata[255:0];
  assign tg6_0_axi_arvalid = m0_arvalid & m0_arready;
  assign tg6_0_axi_arid = m0_arid;
  assign tg6_0_axi_awaddr = {m0_awaddr[31:7], 5'b0};
  assign m0_rdata[1023:768] = tg6_0_axi_rdata;
  assign tg6_0_axi_arburst = m0_arburst;
  assign tg6_0_axi_arsize = m0_arsize;
  assign tg6_0_axi_bready = m0_bready;
  assign tg6_0_axi_wlast = m0_wlast;
  assign tg6_0_axi_awid = m0_awid;
  assign tg6_0_axi_awsize = m0_awsize;
  assign tg6_0_axi_awvalid = m0_awvalid & m0_awready;
  assign tg6_0_axi_aruser = 1'b0;

  //-- port 1
  assign tg0_1_axi_awburst = m1_awburst;
  assign tg0_1_axi_awuser = 1'b0;
  assign tg0_1_axi_arlen = m1_arlen;
  assign tg0_1_axi_arqos = 4'b0;
  assign tg0_1_axi_wstrb = m1_wstrb[31:0];
  assign m1_wready = tg0_1_axi_wready & tg2_1_axi_wready & tg4_1_axi_wready & tg6_1_axi_wready;
  assign m1_rid = tg0_1_axi_rid;
  assign tg0_1_axi_awlen = m1_awlen;
  assign tg0_1_axi_awqos = 4'b0;
  assign tg0_1_axi_wvalid = m1_wvalid & m1_wready;
  assign tg0_1_axi_araddr = {m1_araddr[31:7], 5'b0};
  assign tg0_1_axi_arprot = 3'b0;
  assign tg0_1_axi_awprot = 3'b0;
  assign tg0_1_axi_wdata = m1_wdata[255:0];
  assign tg0_1_axi_arvalid = m1_arvalid & m1_arready;
  assign tg0_1_axi_arid = m1_arid;
  assign tg0_1_axi_awaddr = {m1_awaddr[31:7], 5'b0};
  assign m1_arready = tg0_1_axi_arready & tg2_1_axi_arready & tg4_1_axi_arready & tg6_1_axi_arready;
  assign m1_rdata[255:0] = tg0_1_axi_rdata;
  assign m1_awready = tg0_1_axi_awready & tg2_1_axi_awready & tg4_1_axi_awready & tg6_1_axi_awready;
  assign tg0_1_axi_arburst = m1_arburst;
  assign tg0_1_axi_arsize = m1_arsize;
  assign tg0_1_axi_bready = m1_bready;
  assign m1_rlast = tg0_1_axi_rlast;
  assign tg0_1_axi_wlast = m1_wlast;
  assign tg0_1_axi_awid = m1_awid;
  assign m1_bid = tg0_1_axi_bid;
  assign m1_bvalid = tg0_1_axi_bvalid;
  assign tg0_1_axi_awsize = m1_awsize;
  assign tg0_1_axi_awvalid = m1_awvalid & m1_awready;
  assign tg0_1_axi_aruser = 1'b0;
  assign m1_rvalid = tg0_1_axi_rvalid & tg2_1_axi_rvalid & tg4_1_axi_rvalid & tg6_1_axi_rvalid;

  assign tg2_1_axi_awburst = m1_awburst;
  assign tg2_1_axi_awuser = 1'b0;
  assign tg2_1_axi_arlen = m1_arlen;
  assign tg2_1_axi_arqos = 4'b0;
  assign tg2_1_axi_wstrb = m1_wstrb[63:32];
  assign tg2_1_axi_awlen = m1_awlen;
  assign tg2_1_axi_awqos = 4'b0;
  assign tg2_1_axi_wvalid = m1_wvalid & m1_wready;
  assign tg2_1_axi_araddr = {m1_araddr[31:7], 5'b0};
  assign tg2_1_axi_arprot = 3'b0;
  assign tg2_1_axi_awprot = 3'b0;
  assign tg2_1_axi_wdata = m1_wdata[255:0];
  assign tg2_1_axi_arvalid = m1_arvalid & m1_arready;
  assign tg2_1_axi_arid = m1_arid;
  assign tg2_1_axi_awaddr = {m1_awaddr[31:7], 5'b0};
  assign m1_rdata[511:256] = tg2_1_axi_rdata;
  assign tg2_1_axi_arburst = m1_arburst;
  assign tg2_1_axi_arsize = m1_arsize;
  assign tg2_1_axi_bready = m1_bready;
  assign tg2_1_axi_wlast = m1_wlast;
  assign tg2_1_axi_awid = m1_awid;
  assign tg2_1_axi_awsize = m1_awsize;
  assign tg2_1_axi_awvalid = m1_awvalid & m1_awready;
  assign tg2_1_axi_aruser = 1'b0;

  assign tg4_1_axi_awburst = m1_awburst;
  assign tg4_1_axi_awuser = 1'b0;
  assign tg4_1_axi_arlen = m1_arlen;
  assign tg4_1_axi_arqos = 4'b0;
  assign tg4_1_axi_wstrb = m1_wstrb[95:64];
  assign tg4_1_axi_awlen = m1_awlen;
  assign tg4_1_axi_awqos = 4'b0;
  assign tg4_1_axi_wvalid = m1_wvalid & m1_wready;
  assign tg4_1_axi_araddr = {m1_araddr[31:7], 5'b0};
  assign tg4_1_axi_arprot = 3'b0;
  assign tg4_1_axi_awprot = 3'b0;
  assign tg4_1_axi_wdata = m1_wdata[255:0];
  assign tg4_1_axi_arvalid = m1_arvalid & m1_arready;
  assign tg4_1_axi_arid = m1_arid;
  assign tg4_1_axi_awaddr = {m1_awaddr[31:7], 5'b0};
  assign m1_rdata[767:512] = tg4_1_axi_rdata;
  assign tg4_1_axi_arburst = m1_arburst;
  assign tg4_1_axi_arsize = m1_arsize;
  assign tg4_1_axi_bready = m1_bready;
  assign tg4_1_axi_wlast = m1_wlast;
  assign tg4_1_axi_awid = m1_awid;
  assign tg4_1_axi_awsize = m1_awsize;
  assign tg4_1_axi_awvalid = m1_awvalid & m1_awready;
  assign tg4_1_axi_aruser = 1'b0;

  assign tg6_1_axi_awburst = m1_awburst;
  assign tg6_1_axi_awuser = 1'b0;
  assign tg6_1_axi_arlen = m1_arlen;
  assign tg6_1_axi_arqos = 4'b0;
  assign tg6_1_axi_wstrb = m1_wstrb[127:96];
  assign tg6_1_axi_awlen = m1_awlen;
  assign tg6_1_axi_awqos = 4'b0;
  assign tg6_1_axi_wvalid = m1_wvalid & m1_wready;
  assign tg6_1_axi_araddr = {m1_araddr[31:7], 5'b0};
  assign tg6_1_axi_arprot = 3'b0;
  assign tg6_1_axi_awprot = 3'b0;
  assign tg6_1_axi_wdata = m1_wdata[255:0];
  assign tg6_1_axi_arvalid = m1_arvalid & m1_arready;
  assign tg6_1_axi_arid = m1_arid;
  assign tg6_1_axi_awaddr = {m1_awaddr[31:7], 5'b0};
  assign m1_rdata[1023:768] = tg6_1_axi_rdata;
  assign tg6_1_axi_arburst = m1_arburst;
  assign tg6_1_axi_arsize = m1_arsize;
  assign tg6_1_axi_bready = m1_bready;
  assign tg6_1_axi_wlast = m1_wlast;
  assign tg6_1_axi_awid = m1_awid;
  assign tg6_1_axi_awsize = m1_awsize;
  assign tg6_1_axi_awvalid = m1_awvalid & m1_awready;
  assign tg6_1_axi_aruser = 1'b0;

  //-- port 2
  assign tg1_0_axi_awburst = m2_awburst;
  assign tg1_0_axi_awuser = 1'b0;
  assign tg1_0_axi_arlen = m2_arlen;
  assign tg1_0_axi_arqos = 4'b0;
  assign tg1_0_axi_wstrb = m2_wstrb[31:0];
  assign m2_wready = tg1_0_axi_wready & tg3_0_axi_wready & tg5_0_axi_wready & tg7_0_axi_wready;
  assign m2_rid = tg1_0_axi_rid;
  assign tg1_0_axi_awlen = m2_awlen;
  assign tg1_0_axi_awqos = 4'b0;
  assign tg1_0_axi_wvalid = m2_wvalid & m2_wready;
  assign tg1_0_axi_araddr = {m2_araddr[31:7], 5'b0};
  assign tg1_0_axi_arprot = 3'b0;
  assign tg1_0_axi_awprot = 3'b0;
  assign tg1_0_axi_wdata = m2_wdata[255:0];
  assign tg1_0_axi_arvalid = m2_arvalid & m2_arready;
  assign tg1_0_axi_arid = m2_arid;
  assign tg1_0_axi_awaddr = {m2_awaddr[31:7], 5'b0};
  assign m2_arready = tg1_0_axi_arready & tg3_0_axi_arready & tg5_0_axi_arready & tg7_0_axi_arready;
  assign m2_rdata[255:0] = tg1_0_axi_rdata;
  assign m2_awready = tg1_0_axi_awready & tg3_0_axi_awready & tg5_0_axi_awready & tg7_0_axi_awready;
  assign tg1_0_axi_arburst = m2_arburst;
  assign tg1_0_axi_arsize = m2_arsize;
  assign tg1_0_axi_bready = m2_bready;
  assign m2_rlast = tg1_0_axi_rlast;
  assign tg1_0_axi_wlast = m2_wlast;
  assign tg1_0_axi_awid = m2_awid;
  assign m2_bid = tg1_0_axi_bid;
  assign m2_bvalid = tg1_0_axi_bvalid;
  assign tg1_0_axi_awsize = m2_awsize;
  assign tg1_0_axi_awvalid = m2_awvalid & m2_awready;
  assign tg1_0_axi_aruser = 1'b0;
  assign m2_rvalid = tg1_0_axi_rvalid & tg3_0_axi_rvalid & tg5_0_axi_rvalid & tg7_0_axi_rvalid;

  assign tg3_0_axi_awburst = m2_awburst;
  assign tg3_0_axi_awuser = 1'b0;
  assign tg3_0_axi_arlen = m2_arlen;
  assign tg3_0_axi_arqos = 4'b0;
  assign tg3_0_axi_wstrb = m2_wstrb[63:32];
  assign tg3_0_axi_awlen = m2_awlen;
  assign tg3_0_axi_awqos = 4'b0;
  assign tg3_0_axi_wvalid = m2_wvalid & m2_wready;
  assign tg3_0_axi_araddr = {m2_araddr[31:7], 5'b0};
  assign tg3_0_axi_arprot = 3'b0;
  assign tg3_0_axi_awprot = 3'b0;
  assign tg3_0_axi_wdata = m2_wdata[255:0];
  assign tg3_0_axi_arvalid = m2_arvalid & m2_arready;
  assign tg3_0_axi_arid = m2_arid;
  assign tg3_0_axi_awaddr = {m2_awaddr[31:7], 5'b0};
  assign m2_rdata[511:256] = tg3_0_axi_rdata;
  assign tg3_0_axi_arburst = m2_arburst;
  assign tg3_0_axi_arsize = m2_arsize;
  assign tg3_0_axi_bready = m2_bready;
  assign tg3_0_axi_wlast = m2_wlast;
  assign tg3_0_axi_awid = m2_awid;
  assign tg3_0_axi_awsize = m2_awsize;
  assign tg3_0_axi_awvalid = m2_awvalid & m2_awready;
  assign tg3_0_axi_aruser = 1'b0;

  assign tg5_0_axi_awburst = m2_awburst;
  assign tg5_0_axi_awuser = 1'b0;
  assign tg5_0_axi_arlen = m2_arlen;
  assign tg5_0_axi_arqos = 4'b0;
  assign tg5_0_axi_wstrb = m2_wstrb[95:64];
  assign tg5_0_axi_awlen = m2_awlen;
  assign tg5_0_axi_awqos = 4'b0;
  assign tg5_0_axi_wvalid = m2_wvalid & m2_wready;
  assign tg5_0_axi_araddr = {m2_araddr[31:7], 5'b0};
  assign tg5_0_axi_arprot = 3'b0;
  assign tg5_0_axi_awprot = 3'b0;
  assign tg5_0_axi_wdata = m2_wdata[255:0];
  assign tg5_0_axi_arvalid = m2_arvalid & m2_arready;
  assign tg5_0_axi_arid = m2_arid;
  assign tg5_0_axi_awaddr = {m2_awaddr[31:7], 5'b0};
  assign m2_rdata[767:512] = tg5_0_axi_rdata;
  assign tg5_0_axi_arburst = m2_arburst;
  assign tg5_0_axi_arsize = m2_arsize;
  assign tg5_0_axi_bready = m2_bready;
  assign tg5_0_axi_wlast = m2_wlast;
  assign tg5_0_axi_awid = m2_awid;
  assign tg5_0_axi_awsize = m2_awsize;
  assign tg5_0_axi_awvalid = m2_awvalid & m2_awready;
  assign tg5_0_axi_aruser = 1'b0;

  assign tg7_0_axi_awburst = m2_awburst;
  assign tg7_0_axi_awuser = 1'b0;
  assign tg7_0_axi_arlen = m2_arlen;
  assign tg7_0_axi_arqos = 4'b0;
  assign tg7_0_axi_wstrb = m2_wstrb[127:96];
  assign tg7_0_axi_awlen = m2_awlen;
  assign tg7_0_axi_awqos = 4'b0;
  assign tg7_0_axi_wvalid = m2_wvalid & m2_wready;
  assign tg7_0_axi_araddr = {m2_araddr[31:7], 5'b0};
  assign tg7_0_axi_arprot = 3'b0;
  assign tg7_0_axi_awprot = 3'b0;
  assign tg7_0_axi_wdata = m2_wdata[255:0];
  assign tg7_0_axi_arvalid = m2_arvalid & m2_arready;
  assign tg7_0_axi_arid = m2_arid;
  assign tg7_0_axi_awaddr = {m2_awaddr[31:7], 5'b0};
  assign m2_rdata[1023:768] = tg7_0_axi_rdata;
  assign tg7_0_axi_arburst = m2_arburst;
  assign tg7_0_axi_arsize = m2_arsize;
  assign tg7_0_axi_bready = m2_bready;
  assign tg7_0_axi_wlast = m2_wlast;
  assign tg7_0_axi_awid = m2_awid;
  assign tg7_0_axi_awsize = m2_awsize;
  assign tg7_0_axi_awvalid = m2_awvalid & m2_awready;
  assign tg7_0_axi_aruser = 1'b0;

  //-- port 3
  assign tg1_1_axi_awburst = m3_awburst;
  assign tg1_1_axi_awuser = 1'b0;
  assign tg1_1_axi_arlen = m3_arlen;
  assign tg1_1_axi_arqos = 4'b0;
  assign tg1_1_axi_wstrb = m3_wstrb[31:0];
  assign m3_wready = tg1_1_axi_wready & tg3_1_axi_wready & tg5_1_axi_wready & tg7_1_axi_wready;
  assign m3_rid = tg1_1_axi_rid;
  assign tg1_1_axi_awlen = m3_awlen;
  assign tg1_1_axi_awqos = 4'b0;
  assign tg1_1_axi_wvalid = m3_wvalid & m3_wready;
  assign tg1_1_axi_araddr = {m3_araddr[31:7], 5'b0};
  assign tg1_1_axi_arprot = 3'b0;
  assign tg1_1_axi_awprot = 3'b0;
  assign tg1_1_axi_wdata = m3_wdata[255:0];
  assign tg1_1_axi_arvalid = m3_arvalid & m3_arready;
  assign tg1_1_axi_arid = m3_arid;
  assign tg1_1_axi_awaddr = {m3_awaddr[31:7], 5'b0};
  assign m3_arready = tg1_1_axi_arready & tg3_1_axi_arready & tg5_1_axi_arready & tg7_1_axi_arready;
  assign m3_rdata[255:0] = tg1_1_axi_rdata;
  assign m3_awready = tg1_1_axi_awready & tg3_1_axi_awready & tg5_1_axi_awready & tg7_1_axi_awready;
  assign tg1_1_axi_arburst = m3_arburst;
  assign tg1_1_axi_arsize = m3_arsize;
  assign tg1_1_axi_bready = m3_bready;
  assign m3_rlast = tg1_1_axi_rlast;
  assign tg1_1_axi_wlast = m3_wlast;
  assign tg1_1_axi_awid = m3_awid;
  assign m3_bid = tg1_1_axi_bid;
  assign m3_bvalid = tg1_1_axi_bvalid;
  assign tg1_1_axi_awsize = m3_awsize;
  assign tg1_1_axi_awvalid = m3_awvalid & m3_awready;
  assign tg1_1_axi_aruser = 1'b0;
  assign m3_rvalid = tg1_1_axi_rvalid & tg3_1_axi_rvalid & tg5_1_axi_rvalid & tg7_1_axi_rvalid;

  assign tg3_1_axi_awburst = m3_awburst;
  assign tg3_1_axi_awuser = 1'b0;
  assign tg3_1_axi_arlen = m3_arlen;
  assign tg3_1_axi_arqos = 4'b0;
  assign tg3_1_axi_wstrb = m3_wstrb[63:32];
  assign tg3_1_axi_awlen = m3_awlen;
  assign tg3_1_axi_awqos = 4'b0;
  assign tg3_1_axi_wvalid = m3_wvalid & m3_wready;
  assign tg3_1_axi_araddr = {m3_araddr[31:7], 5'b0};
  assign tg3_1_axi_arprot = 3'b0;
  assign tg3_1_axi_awprot = 3'b0;
  assign tg3_1_axi_wdata = m3_wdata[255:0];
  assign tg3_1_axi_arvalid = m3_arvalid & m3_arready;
  assign tg3_1_axi_arid = m3_arid;
  assign tg3_1_axi_awaddr = {m3_awaddr[31:7], 5'b0};
  assign m3_rdata[511:256] = tg3_1_axi_rdata;
  assign tg3_1_axi_arburst = m3_arburst;
  assign tg3_1_axi_arsize = m3_arsize;
  assign tg3_1_axi_bready = m3_bready;
  assign tg3_1_axi_wlast = m3_wlast;
  assign tg3_1_axi_awid = m3_awid;
  assign tg3_1_axi_awsize = m3_awsize;
  assign tg3_1_axi_awvalid = m3_awvalid & m3_awready;
  assign tg3_1_axi_aruser = 1'b0;

  assign tg5_1_axi_awburst = m3_awburst;
  assign tg5_1_axi_awuser = 1'b0;
  assign tg5_1_axi_arlen = m3_arlen;
  assign tg5_1_axi_arqos = 4'b0;
  assign tg5_1_axi_wstrb = m3_wstrb[95:64];
  assign tg5_1_axi_awlen = m3_awlen;
  assign tg5_1_axi_awqos = 4'b0;
  assign tg5_1_axi_wvalid = m3_wvalid & m3_wready;
  assign tg5_1_axi_araddr = {m3_araddr[31:7], 5'b0};
  assign tg5_1_axi_arprot = 3'b0;
  assign tg5_1_axi_awprot = 3'b0;
  assign tg5_1_axi_wdata = m3_wdata[255:0];
  assign tg5_1_axi_arvalid = m3_arvalid & m3_arready;
  assign tg5_1_axi_arid = m3_arid;
  assign tg5_1_axi_awaddr = {m3_awaddr[31:7], 5'b0};
  assign m3_rdata[767:512] = tg5_1_axi_rdata;
  assign tg5_1_axi_arburst = m3_arburst;
  assign tg5_1_axi_arsize = m3_arsize;
  assign tg5_1_axi_bready = m3_bready;
  assign tg5_1_axi_wlast = m3_wlast;
  assign tg5_1_axi_awid = m3_awid;
  assign tg5_1_axi_awsize = m3_awsize;
  assign tg5_1_axi_awvalid = m3_awvalid & m3_awready;
  assign tg5_1_axi_aruser = 1'b0;

  assign tg7_1_axi_awburst = m3_awburst;
  assign tg7_1_axi_awuser = 1'b0;
  assign tg7_1_axi_arlen = m3_arlen;
  assign tg7_1_axi_arqos = 4'b0;
  assign tg7_1_axi_wstrb = m3_wstrb[127:96];
  assign tg7_1_axi_awlen = m3_awlen;
  assign tg7_1_axi_awqos = 4'b0;
  assign tg7_1_axi_wvalid = m3_wvalid & m3_wready;
  assign tg7_1_axi_araddr = {m3_araddr[31:7], 5'b0};
  assign tg7_1_axi_arprot = 3'b0;
  assign tg7_1_axi_awprot = 3'b0;
  assign tg7_1_axi_wdata = m3_wdata[255:0];
  assign tg7_1_axi_arvalid = m3_arvalid & m3_arready;
  assign tg7_1_axi_arid = m3_arid;
  assign tg7_1_axi_awaddr = {m3_awaddr[31:7], 5'b0};
  assign m3_rdata[1023:768] = tg7_1_axi_rdata;
  assign tg7_1_axi_arburst = m3_arburst;
  assign tg7_1_axi_arsize = m3_arsize;
  assign tg7_1_axi_bready = m3_bready;
  assign tg7_1_axi_wlast = m3_wlast;
  assign tg7_1_axi_awid = m3_awid;
  assign tg7_1_axi_awsize = m3_awsize;
  assign tg7_1_axi_awvalid = m3_awvalid & m3_awready;
  assign tg7_1_axi_aruser = 1'b0;

endmodule
