sim/fir/FGPU_definitions.vhd